// mlp_weights.vh — Placeholder for H=16 (awaiting Colab training)
// Network: 3 -> 16 -> 16 -> 3 SIREN
// Total parameters: 387
// NOTE: These are zero weights — replace with trained weights

initial begin
    weight_mem[  0] = 32'sh00000000;  // L0 w[0][0]
    weight_mem[  1] = 32'sh00000000;  // L0 w[0][1]
    weight_mem[  2] = 32'sh00000000;  // L0 w[0][2]
    weight_mem[  3] = 32'sh00000000;  // L0 w[1][0]
    weight_mem[  4] = 32'sh00000000;  // L0 w[1][1]
    weight_mem[  5] = 32'sh00000000;  // L0 w[1][2]
    weight_mem[  6] = 32'sh00000000;  // L0 w[2][0]
    weight_mem[  7] = 32'sh00000000;  // L0 w[2][1]
    weight_mem[  8] = 32'sh00000000;  // L0 w[2][2]
    weight_mem[  9] = 32'sh00000000;  // L0 w[3][0]
    weight_mem[ 10] = 32'sh00000000;  // L0 w[3][1]
    weight_mem[ 11] = 32'sh00000000;  // L0 w[3][2]
    weight_mem[ 12] = 32'sh00000000;  // L0 w[4][0]
    weight_mem[ 13] = 32'sh00000000;  // L0 w[4][1]
    weight_mem[ 14] = 32'sh00000000;  // L0 w[4][2]
    weight_mem[ 15] = 32'sh00000000;  // L0 w[5][0]
    weight_mem[ 16] = 32'sh00000000;  // L0 w[5][1]
    weight_mem[ 17] = 32'sh00000000;  // L0 w[5][2]
    weight_mem[ 18] = 32'sh00000000;  // L0 w[6][0]
    weight_mem[ 19] = 32'sh00000000;  // L0 w[6][1]
    weight_mem[ 20] = 32'sh00000000;  // L0 w[6][2]
    weight_mem[ 21] = 32'sh00000000;  // L0 w[7][0]
    weight_mem[ 22] = 32'sh00000000;  // L0 w[7][1]
    weight_mem[ 23] = 32'sh00000000;  // L0 w[7][2]
    weight_mem[ 24] = 32'sh00000000;  // L0 w[8][0]
    weight_mem[ 25] = 32'sh00000000;  // L0 w[8][1]
    weight_mem[ 26] = 32'sh00000000;  // L0 w[8][2]
    weight_mem[ 27] = 32'sh00000000;  // L0 w[9][0]
    weight_mem[ 28] = 32'sh00000000;  // L0 w[9][1]
    weight_mem[ 29] = 32'sh00000000;  // L0 w[9][2]
    weight_mem[ 30] = 32'sh00000000;  // L0 w[10][0]
    weight_mem[ 31] = 32'sh00000000;  // L0 w[10][1]
    weight_mem[ 32] = 32'sh00000000;  // L0 w[10][2]
    weight_mem[ 33] = 32'sh00000000;  // L0 w[11][0]
    weight_mem[ 34] = 32'sh00000000;  // L0 w[11][1]
    weight_mem[ 35] = 32'sh00000000;  // L0 w[11][2]
    weight_mem[ 36] = 32'sh00000000;  // L0 w[12][0]
    weight_mem[ 37] = 32'sh00000000;  // L0 w[12][1]
    weight_mem[ 38] = 32'sh00000000;  // L0 w[12][2]
    weight_mem[ 39] = 32'sh00000000;  // L0 w[13][0]
    weight_mem[ 40] = 32'sh00000000;  // L0 w[13][1]
    weight_mem[ 41] = 32'sh00000000;  // L0 w[13][2]
    weight_mem[ 42] = 32'sh00000000;  // L0 w[14][0]
    weight_mem[ 43] = 32'sh00000000;  // L0 w[14][1]
    weight_mem[ 44] = 32'sh00000000;  // L0 w[14][2]
    weight_mem[ 45] = 32'sh00000000;  // L0 w[15][0]
    weight_mem[ 46] = 32'sh00000000;  // L0 w[15][1]
    weight_mem[ 47] = 32'sh00000000;  // L0 w[15][2]
    weight_mem[ 48] = 32'sh00000000;  // L0 b[0]
    weight_mem[ 49] = 32'sh00000000;  // L0 b[1]
    weight_mem[ 50] = 32'sh00000000;  // L0 b[2]
    weight_mem[ 51] = 32'sh00000000;  // L0 b[3]
    weight_mem[ 52] = 32'sh00000000;  // L0 b[4]
    weight_mem[ 53] = 32'sh00000000;  // L0 b[5]
    weight_mem[ 54] = 32'sh00000000;  // L0 b[6]
    weight_mem[ 55] = 32'sh00000000;  // L0 b[7]
    weight_mem[ 56] = 32'sh00000000;  // L0 b[8]
    weight_mem[ 57] = 32'sh00000000;  // L0 b[9]
    weight_mem[ 58] = 32'sh00000000;  // L0 b[10]
    weight_mem[ 59] = 32'sh00000000;  // L0 b[11]
    weight_mem[ 60] = 32'sh00000000;  // L0 b[12]
    weight_mem[ 61] = 32'sh00000000;  // L0 b[13]
    weight_mem[ 62] = 32'sh00000000;  // L0 b[14]
    weight_mem[ 63] = 32'sh00000000;  // L0 b[15]
    weight_mem[ 64] = 32'sh00000000;  // L1 w[0][0]
    weight_mem[ 65] = 32'sh00000000;  // L1 w[0][1]
    weight_mem[ 66] = 32'sh00000000;  // L1 w[0][2]
    weight_mem[ 67] = 32'sh00000000;  // L1 w[0][3]
    weight_mem[ 68] = 32'sh00000000;  // L1 w[0][4]
    weight_mem[ 69] = 32'sh00000000;  // L1 w[0][5]
    weight_mem[ 70] = 32'sh00000000;  // L1 w[0][6]
    weight_mem[ 71] = 32'sh00000000;  // L1 w[0][7]
    weight_mem[ 72] = 32'sh00000000;  // L1 w[0][8]
    weight_mem[ 73] = 32'sh00000000;  // L1 w[0][9]
    weight_mem[ 74] = 32'sh00000000;  // L1 w[0][10]
    weight_mem[ 75] = 32'sh00000000;  // L1 w[0][11]
    weight_mem[ 76] = 32'sh00000000;  // L1 w[0][12]
    weight_mem[ 77] = 32'sh00000000;  // L1 w[0][13]
    weight_mem[ 78] = 32'sh00000000;  // L1 w[0][14]
    weight_mem[ 79] = 32'sh00000000;  // L1 w[0][15]
    weight_mem[ 80] = 32'sh00000000;  // L1 w[1][0]
    weight_mem[ 81] = 32'sh00000000;  // L1 w[1][1]
    weight_mem[ 82] = 32'sh00000000;  // L1 w[1][2]
    weight_mem[ 83] = 32'sh00000000;  // L1 w[1][3]
    weight_mem[ 84] = 32'sh00000000;  // L1 w[1][4]
    weight_mem[ 85] = 32'sh00000000;  // L1 w[1][5]
    weight_mem[ 86] = 32'sh00000000;  // L1 w[1][6]
    weight_mem[ 87] = 32'sh00000000;  // L1 w[1][7]
    weight_mem[ 88] = 32'sh00000000;  // L1 w[1][8]
    weight_mem[ 89] = 32'sh00000000;  // L1 w[1][9]
    weight_mem[ 90] = 32'sh00000000;  // L1 w[1][10]
    weight_mem[ 91] = 32'sh00000000;  // L1 w[1][11]
    weight_mem[ 92] = 32'sh00000000;  // L1 w[1][12]
    weight_mem[ 93] = 32'sh00000000;  // L1 w[1][13]
    weight_mem[ 94] = 32'sh00000000;  // L1 w[1][14]
    weight_mem[ 95] = 32'sh00000000;  // L1 w[1][15]
    weight_mem[ 96] = 32'sh00000000;  // L1 w[2][0]
    weight_mem[ 97] = 32'sh00000000;  // L1 w[2][1]
    weight_mem[ 98] = 32'sh00000000;  // L1 w[2][2]
    weight_mem[ 99] = 32'sh00000000;  // L1 w[2][3]
    weight_mem[100] = 32'sh00000000;  // L1 w[2][4]
    weight_mem[101] = 32'sh00000000;  // L1 w[2][5]
    weight_mem[102] = 32'sh00000000;  // L1 w[2][6]
    weight_mem[103] = 32'sh00000000;  // L1 w[2][7]
    weight_mem[104] = 32'sh00000000;  // L1 w[2][8]
    weight_mem[105] = 32'sh00000000;  // L1 w[2][9]
    weight_mem[106] = 32'sh00000000;  // L1 w[2][10]
    weight_mem[107] = 32'sh00000000;  // L1 w[2][11]
    weight_mem[108] = 32'sh00000000;  // L1 w[2][12]
    weight_mem[109] = 32'sh00000000;  // L1 w[2][13]
    weight_mem[110] = 32'sh00000000;  // L1 w[2][14]
    weight_mem[111] = 32'sh00000000;  // L1 w[2][15]
    weight_mem[112] = 32'sh00000000;  // L1 w[3][0]
    weight_mem[113] = 32'sh00000000;  // L1 w[3][1]
    weight_mem[114] = 32'sh00000000;  // L1 w[3][2]
    weight_mem[115] = 32'sh00000000;  // L1 w[3][3]
    weight_mem[116] = 32'sh00000000;  // L1 w[3][4]
    weight_mem[117] = 32'sh00000000;  // L1 w[3][5]
    weight_mem[118] = 32'sh00000000;  // L1 w[3][6]
    weight_mem[119] = 32'sh00000000;  // L1 w[3][7]
    weight_mem[120] = 32'sh00000000;  // L1 w[3][8]
    weight_mem[121] = 32'sh00000000;  // L1 w[3][9]
    weight_mem[122] = 32'sh00000000;  // L1 w[3][10]
    weight_mem[123] = 32'sh00000000;  // L1 w[3][11]
    weight_mem[124] = 32'sh00000000;  // L1 w[3][12]
    weight_mem[125] = 32'sh00000000;  // L1 w[3][13]
    weight_mem[126] = 32'sh00000000;  // L1 w[3][14]
    weight_mem[127] = 32'sh00000000;  // L1 w[3][15]
    weight_mem[128] = 32'sh00000000;  // L1 w[4][0]
    weight_mem[129] = 32'sh00000000;  // L1 w[4][1]
    weight_mem[130] = 32'sh00000000;  // L1 w[4][2]
    weight_mem[131] = 32'sh00000000;  // L1 w[4][3]
    weight_mem[132] = 32'sh00000000;  // L1 w[4][4]
    weight_mem[133] = 32'sh00000000;  // L1 w[4][5]
    weight_mem[134] = 32'sh00000000;  // L1 w[4][6]
    weight_mem[135] = 32'sh00000000;  // L1 w[4][7]
    weight_mem[136] = 32'sh00000000;  // L1 w[4][8]
    weight_mem[137] = 32'sh00000000;  // L1 w[4][9]
    weight_mem[138] = 32'sh00000000;  // L1 w[4][10]
    weight_mem[139] = 32'sh00000000;  // L1 w[4][11]
    weight_mem[140] = 32'sh00000000;  // L1 w[4][12]
    weight_mem[141] = 32'sh00000000;  // L1 w[4][13]
    weight_mem[142] = 32'sh00000000;  // L1 w[4][14]
    weight_mem[143] = 32'sh00000000;  // L1 w[4][15]
    weight_mem[144] = 32'sh00000000;  // L1 w[5][0]
    weight_mem[145] = 32'sh00000000;  // L1 w[5][1]
    weight_mem[146] = 32'sh00000000;  // L1 w[5][2]
    weight_mem[147] = 32'sh00000000;  // L1 w[5][3]
    weight_mem[148] = 32'sh00000000;  // L1 w[5][4]
    weight_mem[149] = 32'sh00000000;  // L1 w[5][5]
    weight_mem[150] = 32'sh00000000;  // L1 w[5][6]
    weight_mem[151] = 32'sh00000000;  // L1 w[5][7]
    weight_mem[152] = 32'sh00000000;  // L1 w[5][8]
    weight_mem[153] = 32'sh00000000;  // L1 w[5][9]
    weight_mem[154] = 32'sh00000000;  // L1 w[5][10]
    weight_mem[155] = 32'sh00000000;  // L1 w[5][11]
    weight_mem[156] = 32'sh00000000;  // L1 w[5][12]
    weight_mem[157] = 32'sh00000000;  // L1 w[5][13]
    weight_mem[158] = 32'sh00000000;  // L1 w[5][14]
    weight_mem[159] = 32'sh00000000;  // L1 w[5][15]
    weight_mem[160] = 32'sh00000000;  // L1 w[6][0]
    weight_mem[161] = 32'sh00000000;  // L1 w[6][1]
    weight_mem[162] = 32'sh00000000;  // L1 w[6][2]
    weight_mem[163] = 32'sh00000000;  // L1 w[6][3]
    weight_mem[164] = 32'sh00000000;  // L1 w[6][4]
    weight_mem[165] = 32'sh00000000;  // L1 w[6][5]
    weight_mem[166] = 32'sh00000000;  // L1 w[6][6]
    weight_mem[167] = 32'sh00000000;  // L1 w[6][7]
    weight_mem[168] = 32'sh00000000;  // L1 w[6][8]
    weight_mem[169] = 32'sh00000000;  // L1 w[6][9]
    weight_mem[170] = 32'sh00000000;  // L1 w[6][10]
    weight_mem[171] = 32'sh00000000;  // L1 w[6][11]
    weight_mem[172] = 32'sh00000000;  // L1 w[6][12]
    weight_mem[173] = 32'sh00000000;  // L1 w[6][13]
    weight_mem[174] = 32'sh00000000;  // L1 w[6][14]
    weight_mem[175] = 32'sh00000000;  // L1 w[6][15]
    weight_mem[176] = 32'sh00000000;  // L1 w[7][0]
    weight_mem[177] = 32'sh00000000;  // L1 w[7][1]
    weight_mem[178] = 32'sh00000000;  // L1 w[7][2]
    weight_mem[179] = 32'sh00000000;  // L1 w[7][3]
    weight_mem[180] = 32'sh00000000;  // L1 w[7][4]
    weight_mem[181] = 32'sh00000000;  // L1 w[7][5]
    weight_mem[182] = 32'sh00000000;  // L1 w[7][6]
    weight_mem[183] = 32'sh00000000;  // L1 w[7][7]
    weight_mem[184] = 32'sh00000000;  // L1 w[7][8]
    weight_mem[185] = 32'sh00000000;  // L1 w[7][9]
    weight_mem[186] = 32'sh00000000;  // L1 w[7][10]
    weight_mem[187] = 32'sh00000000;  // L1 w[7][11]
    weight_mem[188] = 32'sh00000000;  // L1 w[7][12]
    weight_mem[189] = 32'sh00000000;  // L1 w[7][13]
    weight_mem[190] = 32'sh00000000;  // L1 w[7][14]
    weight_mem[191] = 32'sh00000000;  // L1 w[7][15]
    weight_mem[192] = 32'sh00000000;  // L1 w[8][0]
    weight_mem[193] = 32'sh00000000;  // L1 w[8][1]
    weight_mem[194] = 32'sh00000000;  // L1 w[8][2]
    weight_mem[195] = 32'sh00000000;  // L1 w[8][3]
    weight_mem[196] = 32'sh00000000;  // L1 w[8][4]
    weight_mem[197] = 32'sh00000000;  // L1 w[8][5]
    weight_mem[198] = 32'sh00000000;  // L1 w[8][6]
    weight_mem[199] = 32'sh00000000;  // L1 w[8][7]
    weight_mem[200] = 32'sh00000000;  // L1 w[8][8]
    weight_mem[201] = 32'sh00000000;  // L1 w[8][9]
    weight_mem[202] = 32'sh00000000;  // L1 w[8][10]
    weight_mem[203] = 32'sh00000000;  // L1 w[8][11]
    weight_mem[204] = 32'sh00000000;  // L1 w[8][12]
    weight_mem[205] = 32'sh00000000;  // L1 w[8][13]
    weight_mem[206] = 32'sh00000000;  // L1 w[8][14]
    weight_mem[207] = 32'sh00000000;  // L1 w[8][15]
    weight_mem[208] = 32'sh00000000;  // L1 w[9][0]
    weight_mem[209] = 32'sh00000000;  // L1 w[9][1]
    weight_mem[210] = 32'sh00000000;  // L1 w[9][2]
    weight_mem[211] = 32'sh00000000;  // L1 w[9][3]
    weight_mem[212] = 32'sh00000000;  // L1 w[9][4]
    weight_mem[213] = 32'sh00000000;  // L1 w[9][5]
    weight_mem[214] = 32'sh00000000;  // L1 w[9][6]
    weight_mem[215] = 32'sh00000000;  // L1 w[9][7]
    weight_mem[216] = 32'sh00000000;  // L1 w[9][8]
    weight_mem[217] = 32'sh00000000;  // L1 w[9][9]
    weight_mem[218] = 32'sh00000000;  // L1 w[9][10]
    weight_mem[219] = 32'sh00000000;  // L1 w[9][11]
    weight_mem[220] = 32'sh00000000;  // L1 w[9][12]
    weight_mem[221] = 32'sh00000000;  // L1 w[9][13]
    weight_mem[222] = 32'sh00000000;  // L1 w[9][14]
    weight_mem[223] = 32'sh00000000;  // L1 w[9][15]
    weight_mem[224] = 32'sh00000000;  // L1 w[10][0]
    weight_mem[225] = 32'sh00000000;  // L1 w[10][1]
    weight_mem[226] = 32'sh00000000;  // L1 w[10][2]
    weight_mem[227] = 32'sh00000000;  // L1 w[10][3]
    weight_mem[228] = 32'sh00000000;  // L1 w[10][4]
    weight_mem[229] = 32'sh00000000;  // L1 w[10][5]
    weight_mem[230] = 32'sh00000000;  // L1 w[10][6]
    weight_mem[231] = 32'sh00000000;  // L1 w[10][7]
    weight_mem[232] = 32'sh00000000;  // L1 w[10][8]
    weight_mem[233] = 32'sh00000000;  // L1 w[10][9]
    weight_mem[234] = 32'sh00000000;  // L1 w[10][10]
    weight_mem[235] = 32'sh00000000;  // L1 w[10][11]
    weight_mem[236] = 32'sh00000000;  // L1 w[10][12]
    weight_mem[237] = 32'sh00000000;  // L1 w[10][13]
    weight_mem[238] = 32'sh00000000;  // L1 w[10][14]
    weight_mem[239] = 32'sh00000000;  // L1 w[10][15]
    weight_mem[240] = 32'sh00000000;  // L1 w[11][0]
    weight_mem[241] = 32'sh00000000;  // L1 w[11][1]
    weight_mem[242] = 32'sh00000000;  // L1 w[11][2]
    weight_mem[243] = 32'sh00000000;  // L1 w[11][3]
    weight_mem[244] = 32'sh00000000;  // L1 w[11][4]
    weight_mem[245] = 32'sh00000000;  // L1 w[11][5]
    weight_mem[246] = 32'sh00000000;  // L1 w[11][6]
    weight_mem[247] = 32'sh00000000;  // L1 w[11][7]
    weight_mem[248] = 32'sh00000000;  // L1 w[11][8]
    weight_mem[249] = 32'sh00000000;  // L1 w[11][9]
    weight_mem[250] = 32'sh00000000;  // L1 w[11][10]
    weight_mem[251] = 32'sh00000000;  // L1 w[11][11]
    weight_mem[252] = 32'sh00000000;  // L1 w[11][12]
    weight_mem[253] = 32'sh00000000;  // L1 w[11][13]
    weight_mem[254] = 32'sh00000000;  // L1 w[11][14]
    weight_mem[255] = 32'sh00000000;  // L1 w[11][15]
    weight_mem[256] = 32'sh00000000;  // L1 w[12][0]
    weight_mem[257] = 32'sh00000000;  // L1 w[12][1]
    weight_mem[258] = 32'sh00000000;  // L1 w[12][2]
    weight_mem[259] = 32'sh00000000;  // L1 w[12][3]
    weight_mem[260] = 32'sh00000000;  // L1 w[12][4]
    weight_mem[261] = 32'sh00000000;  // L1 w[12][5]
    weight_mem[262] = 32'sh00000000;  // L1 w[12][6]
    weight_mem[263] = 32'sh00000000;  // L1 w[12][7]
    weight_mem[264] = 32'sh00000000;  // L1 w[12][8]
    weight_mem[265] = 32'sh00000000;  // L1 w[12][9]
    weight_mem[266] = 32'sh00000000;  // L1 w[12][10]
    weight_mem[267] = 32'sh00000000;  // L1 w[12][11]
    weight_mem[268] = 32'sh00000000;  // L1 w[12][12]
    weight_mem[269] = 32'sh00000000;  // L1 w[12][13]
    weight_mem[270] = 32'sh00000000;  // L1 w[12][14]
    weight_mem[271] = 32'sh00000000;  // L1 w[12][15]
    weight_mem[272] = 32'sh00000000;  // L1 w[13][0]
    weight_mem[273] = 32'sh00000000;  // L1 w[13][1]
    weight_mem[274] = 32'sh00000000;  // L1 w[13][2]
    weight_mem[275] = 32'sh00000000;  // L1 w[13][3]
    weight_mem[276] = 32'sh00000000;  // L1 w[13][4]
    weight_mem[277] = 32'sh00000000;  // L1 w[13][5]
    weight_mem[278] = 32'sh00000000;  // L1 w[13][6]
    weight_mem[279] = 32'sh00000000;  // L1 w[13][7]
    weight_mem[280] = 32'sh00000000;  // L1 w[13][8]
    weight_mem[281] = 32'sh00000000;  // L1 w[13][9]
    weight_mem[282] = 32'sh00000000;  // L1 w[13][10]
    weight_mem[283] = 32'sh00000000;  // L1 w[13][11]
    weight_mem[284] = 32'sh00000000;  // L1 w[13][12]
    weight_mem[285] = 32'sh00000000;  // L1 w[13][13]
    weight_mem[286] = 32'sh00000000;  // L1 w[13][14]
    weight_mem[287] = 32'sh00000000;  // L1 w[13][15]
    weight_mem[288] = 32'sh00000000;  // L1 w[14][0]
    weight_mem[289] = 32'sh00000000;  // L1 w[14][1]
    weight_mem[290] = 32'sh00000000;  // L1 w[14][2]
    weight_mem[291] = 32'sh00000000;  // L1 w[14][3]
    weight_mem[292] = 32'sh00000000;  // L1 w[14][4]
    weight_mem[293] = 32'sh00000000;  // L1 w[14][5]
    weight_mem[294] = 32'sh00000000;  // L1 w[14][6]
    weight_mem[295] = 32'sh00000000;  // L1 w[14][7]
    weight_mem[296] = 32'sh00000000;  // L1 w[14][8]
    weight_mem[297] = 32'sh00000000;  // L1 w[14][9]
    weight_mem[298] = 32'sh00000000;  // L1 w[14][10]
    weight_mem[299] = 32'sh00000000;  // L1 w[14][11]
    weight_mem[300] = 32'sh00000000;  // L1 w[14][12]
    weight_mem[301] = 32'sh00000000;  // L1 w[14][13]
    weight_mem[302] = 32'sh00000000;  // L1 w[14][14]
    weight_mem[303] = 32'sh00000000;  // L1 w[14][15]
    weight_mem[304] = 32'sh00000000;  // L1 w[15][0]
    weight_mem[305] = 32'sh00000000;  // L1 w[15][1]
    weight_mem[306] = 32'sh00000000;  // L1 w[15][2]
    weight_mem[307] = 32'sh00000000;  // L1 w[15][3]
    weight_mem[308] = 32'sh00000000;  // L1 w[15][4]
    weight_mem[309] = 32'sh00000000;  // L1 w[15][5]
    weight_mem[310] = 32'sh00000000;  // L1 w[15][6]
    weight_mem[311] = 32'sh00000000;  // L1 w[15][7]
    weight_mem[312] = 32'sh00000000;  // L1 w[15][8]
    weight_mem[313] = 32'sh00000000;  // L1 w[15][9]
    weight_mem[314] = 32'sh00000000;  // L1 w[15][10]
    weight_mem[315] = 32'sh00000000;  // L1 w[15][11]
    weight_mem[316] = 32'sh00000000;  // L1 w[15][12]
    weight_mem[317] = 32'sh00000000;  // L1 w[15][13]
    weight_mem[318] = 32'sh00000000;  // L1 w[15][14]
    weight_mem[319] = 32'sh00000000;  // L1 w[15][15]
    weight_mem[320] = 32'sh00000000;  // L1 b[0]
    weight_mem[321] = 32'sh00000000;  // L1 b[1]
    weight_mem[322] = 32'sh00000000;  // L1 b[2]
    weight_mem[323] = 32'sh00000000;  // L1 b[3]
    weight_mem[324] = 32'sh00000000;  // L1 b[4]
    weight_mem[325] = 32'sh00000000;  // L1 b[5]
    weight_mem[326] = 32'sh00000000;  // L1 b[6]
    weight_mem[327] = 32'sh00000000;  // L1 b[7]
    weight_mem[328] = 32'sh00000000;  // L1 b[8]
    weight_mem[329] = 32'sh00000000;  // L1 b[9]
    weight_mem[330] = 32'sh00000000;  // L1 b[10]
    weight_mem[331] = 32'sh00000000;  // L1 b[11]
    weight_mem[332] = 32'sh00000000;  // L1 b[12]
    weight_mem[333] = 32'sh00000000;  // L1 b[13]
    weight_mem[334] = 32'sh00000000;  // L1 b[14]
    weight_mem[335] = 32'sh00000000;  // L1 b[15]
    weight_mem[336] = 32'sh00000000;  // L2 w[0][0]
    weight_mem[337] = 32'sh00000000;  // L2 w[0][1]
    weight_mem[338] = 32'sh00000000;  // L2 w[0][2]
    weight_mem[339] = 32'sh00000000;  // L2 w[0][3]
    weight_mem[340] = 32'sh00000000;  // L2 w[0][4]
    weight_mem[341] = 32'sh00000000;  // L2 w[0][5]
    weight_mem[342] = 32'sh00000000;  // L2 w[0][6]
    weight_mem[343] = 32'sh00000000;  // L2 w[0][7]
    weight_mem[344] = 32'sh00000000;  // L2 w[0][8]
    weight_mem[345] = 32'sh00000000;  // L2 w[0][9]
    weight_mem[346] = 32'sh00000000;  // L2 w[0][10]
    weight_mem[347] = 32'sh00000000;  // L2 w[0][11]
    weight_mem[348] = 32'sh00000000;  // L2 w[0][12]
    weight_mem[349] = 32'sh00000000;  // L2 w[0][13]
    weight_mem[350] = 32'sh00000000;  // L2 w[0][14]
    weight_mem[351] = 32'sh00000000;  // L2 w[0][15]
    weight_mem[352] = 32'sh00000000;  // L2 w[1][0]
    weight_mem[353] = 32'sh00000000;  // L2 w[1][1]
    weight_mem[354] = 32'sh00000000;  // L2 w[1][2]
    weight_mem[355] = 32'sh00000000;  // L2 w[1][3]
    weight_mem[356] = 32'sh00000000;  // L2 w[1][4]
    weight_mem[357] = 32'sh00000000;  // L2 w[1][5]
    weight_mem[358] = 32'sh00000000;  // L2 w[1][6]
    weight_mem[359] = 32'sh00000000;  // L2 w[1][7]
    weight_mem[360] = 32'sh00000000;  // L2 w[1][8]
    weight_mem[361] = 32'sh00000000;  // L2 w[1][9]
    weight_mem[362] = 32'sh00000000;  // L2 w[1][10]
    weight_mem[363] = 32'sh00000000;  // L2 w[1][11]
    weight_mem[364] = 32'sh00000000;  // L2 w[1][12]
    weight_mem[365] = 32'sh00000000;  // L2 w[1][13]
    weight_mem[366] = 32'sh00000000;  // L2 w[1][14]
    weight_mem[367] = 32'sh00000000;  // L2 w[1][15]
    weight_mem[368] = 32'sh00000000;  // L2 w[2][0]
    weight_mem[369] = 32'sh00000000;  // L2 w[2][1]
    weight_mem[370] = 32'sh00000000;  // L2 w[2][2]
    weight_mem[371] = 32'sh00000000;  // L2 w[2][3]
    weight_mem[372] = 32'sh00000000;  // L2 w[2][4]
    weight_mem[373] = 32'sh00000000;  // L2 w[2][5]
    weight_mem[374] = 32'sh00000000;  // L2 w[2][6]
    weight_mem[375] = 32'sh00000000;  // L2 w[2][7]
    weight_mem[376] = 32'sh00000000;  // L2 w[2][8]
    weight_mem[377] = 32'sh00000000;  // L2 w[2][9]
    weight_mem[378] = 32'sh00000000;  // L2 w[2][10]
    weight_mem[379] = 32'sh00000000;  // L2 w[2][11]
    weight_mem[380] = 32'sh00000000;  // L2 w[2][12]
    weight_mem[381] = 32'sh00000000;  // L2 w[2][13]
    weight_mem[382] = 32'sh00000000;  // L2 w[2][14]
    weight_mem[383] = 32'sh00000000;  // L2 w[2][15]
    weight_mem[384] = 32'sh00000000;  // L2 b[0]
    weight_mem[385] = 32'sh00000000;  // L2 b[1]
    weight_mem[386] = 32'sh00000000;  // L2 b[2]
end
