// mlp_weights.vh — Dual-pattern morph weights
// Pattern A: euler_vorticity 32H
// Pattern B: fracture 32H
// Parameters per pattern: 1283

// Pattern A weights
initial begin
    weight_mem[   0] = 32'shFF09AE81;
    weight_mem[   1] = 32'sh38ACBB80;
    weight_mem[   2] = 32'shD9655200;
    weight_mem[   3] = 32'sh05DC23E0;
    weight_mem[   4] = 32'shEEED9520;
    weight_mem[   5] = 32'shCA5DF700;
    weight_mem[   6] = 32'sh1D738CE0;
    weight_mem[   7] = 32'shD43A0280;
    weight_mem[   8] = 32'sh2A17E640;
    weight_mem[   9] = 32'shF453B160;
    weight_mem[  10] = 32'sh337F8080;
    weight_mem[  11] = 32'sh007CEFE1;
    weight_mem[  12] = 32'shD184F080;
    weight_mem[  13] = 32'shEF752600;
    weight_mem[  14] = 32'sh38FAD4C0;
    weight_mem[  15] = 32'sh34C47E00;
    weight_mem[  16] = 32'shEBBFF740;
    weight_mem[  17] = 32'sh32526E00;
    weight_mem[  18] = 32'sh01DF4D3C;
    weight_mem[  19] = 32'sh057025D0;
    weight_mem[  20] = 32'shF7EE4650;
    weight_mem[  21] = 32'shEC1193E0;
    weight_mem[  22] = 32'sh01B86D42;
    weight_mem[  23] = 32'shFEBDC0E0;
    weight_mem[  24] = 32'shC8C8A580;
    weight_mem[  25] = 32'shF3F41040;
    weight_mem[  26] = 32'sh3491A840;
    weight_mem[  27] = 32'shFFBBEEEA;
    weight_mem[  28] = 32'shC5996280;
    weight_mem[  29] = 32'sh176C38C0;
    weight_mem[  30] = 32'sh096D45E0;
    weight_mem[  31] = 32'shC8337CC0;
    weight_mem[  32] = 32'sh26F01480;
    weight_mem[  33] = 32'shCDE32C00;
    weight_mem[  34] = 32'shE395FAC0;
    weight_mem[  35] = 32'sh053B8960;
    weight_mem[  36] = 32'sh2B7BAA00;
    weight_mem[  37] = 32'sh12699E80;
    weight_mem[  38] = 32'sh25F37400;
    weight_mem[  39] = 32'sh011474F2;
    weight_mem[  40] = 32'shC861D680;
    weight_mem[  41] = 32'shE8B06B80;
    weight_mem[  42] = 32'sh01136156;
    weight_mem[  43] = 32'shC7F7CD00;
    weight_mem[  44] = 32'sh27219000;
    weight_mem[  45] = 32'shE869F4C0;
    weight_mem[  46] = 32'shB2037380;
    weight_mem[  47] = 32'shCC7A3840;
    weight_mem[  48] = 32'shC8A26F80;
    weight_mem[  49] = 32'shF5B2EAD0;
    weight_mem[  50] = 32'sh31C23500;
    weight_mem[  51] = 32'shFD725070;
    weight_mem[  52] = 32'sh02FBB304;
    weight_mem[  53] = 32'shFAF3ACC0;
    weight_mem[  54] = 32'sh2BADBE80;
    weight_mem[  55] = 32'sh09543770;
    weight_mem[  56] = 32'sh1B44E260;
    weight_mem[  57] = 32'sh33BE0380;
    weight_mem[  58] = 32'shECF797E0;
    weight_mem[  59] = 32'sh32B23B80;
    weight_mem[  60] = 32'shCEA3ED00;
    weight_mem[  61] = 32'sh0AB881D0;
    weight_mem[  62] = 32'shFD5AFF88;
    weight_mem[  63] = 32'shC48888C0;
    weight_mem[  64] = 32'sh0E198B60;
    weight_mem[  65] = 32'sh005CE2B2;
    weight_mem[  66] = 32'shF5B5ED90;
    weight_mem[  67] = 32'sh05E60FF8;
    weight_mem[  68] = 32'sh139F63E0;
    weight_mem[  69] = 32'shD2E34980;
    weight_mem[  70] = 32'shF19707D0;
    weight_mem[  71] = 32'shDF877EC0;
    weight_mem[  72] = 32'sh0028C648;
    weight_mem[  73] = 32'shC558E400;
    weight_mem[  74] = 32'sh19661C40;
    weight_mem[  75] = 32'shFB482020;
    weight_mem[  76] = 32'sh384AE580;
    weight_mem[  77] = 32'shD3DF4700;
    weight_mem[  78] = 32'sh0CE60520;
    weight_mem[  79] = 32'sh1FFF0CC0;
    weight_mem[  80] = 32'sh05B8A2C0;
    weight_mem[  81] = 32'sh2664ECC0;
    weight_mem[  82] = 32'sh2D6060C0;
    weight_mem[  83] = 32'sh01491C38;
    weight_mem[  84] = 32'shFF8A6507;
    weight_mem[  85] = 32'shC5B0EA40;
    weight_mem[  86] = 32'sh214A3340;
    weight_mem[  87] = 32'shF768E5E0;
    weight_mem[  88] = 32'sh29819D80;
    weight_mem[  89] = 32'sh1D310200;
    weight_mem[  90] = 32'shFFD9031E;
    weight_mem[  91] = 32'shC5E0CF80;
    weight_mem[  92] = 32'sh1E4A1000;
    weight_mem[  93] = 32'sh269C4000;
    weight_mem[  94] = 32'shF4C23420;
    weight_mem[  95] = 32'shDE345B80;
    weight_mem[  96] = 32'sh57FFD480;
    weight_mem[  97] = 32'shE6BC0780;
    weight_mem[  98] = 32'sh2C30DCC0;
    weight_mem[  99] = 32'shE3AC38E0;
    weight_mem[ 100] = 32'sh37E2D900;
    weight_mem[ 101] = 32'sh60F6BE80;
    weight_mem[ 102] = 32'sh4129F380;
    weight_mem[ 103] = 32'shBA562580;
    weight_mem[ 104] = 32'shB9901B00;
    weight_mem[ 105] = 32'sh2D391380;
    weight_mem[ 106] = 32'sh0A709060;
    weight_mem[ 107] = 32'sh30205F00;
    weight_mem[ 108] = 32'shAA7C3E80;
    weight_mem[ 109] = 32'sh36B372C0;
    weight_mem[ 110] = 32'sh0986A590;
    weight_mem[ 111] = 32'sh0D0BF7F0;
    weight_mem[ 112] = 32'shC8509780;
    weight_mem[ 113] = 32'shCD2E1880;
    weight_mem[ 114] = 32'shE55E2440;
    weight_mem[ 115] = 32'sh5EBDF280;
    weight_mem[ 116] = 32'sh2614F380;
    weight_mem[ 117] = 32'shB3065480;
    weight_mem[ 118] = 32'shE27F1540;
    weight_mem[ 119] = 32'shA0F43380;
    weight_mem[ 120] = 32'sh22636100;
    weight_mem[ 121] = 32'sh43C12380;
    weight_mem[ 122] = 32'shC2E84080;
    weight_mem[ 123] = 32'sh118E8B60;
    weight_mem[ 124] = 32'sh29B17F00;
    weight_mem[ 125] = 32'shDA544A80;
    weight_mem[ 126] = 32'shD5173C40;
    weight_mem[ 127] = 32'sh1B007A40;
    weight_mem[ 128] = 32'shF966EA48;
    weight_mem[ 129] = 32'sh0190AC12;
    weight_mem[ 130] = 32'shFE2F8A88;
    weight_mem[ 131] = 32'sh03707194;
    weight_mem[ 132] = 32'shFFD21B8E;
    weight_mem[ 133] = 32'sh053633F0;
    weight_mem[ 134] = 32'shFFD56C54;
    weight_mem[ 135] = 32'shFB2EE4B8;
    weight_mem[ 136] = 32'sh01C217F0;
    weight_mem[ 137] = 32'sh014B0D62;
    weight_mem[ 138] = 32'sh017D1022;
    weight_mem[ 139] = 32'sh035D6A84;
    weight_mem[ 140] = 32'sh0111890A;
    weight_mem[ 141] = 32'sh02315388;
    weight_mem[ 142] = 32'shFBF5E938;
    weight_mem[ 143] = 32'sh0194DEA0;
    weight_mem[ 144] = 32'shFE35A11A;
    weight_mem[ 145] = 32'sh04383648;
    weight_mem[ 146] = 32'shFEB673E2;
    weight_mem[ 147] = 32'shFC045F1C;
    weight_mem[ 148] = 32'shFC84FC4C;
    weight_mem[ 149] = 32'sh0152AA52;
    weight_mem[ 150] = 32'shFECF6E1C;
    weight_mem[ 151] = 32'shFF5EB321;
    weight_mem[ 152] = 32'shFC0FDED8;
    weight_mem[ 153] = 32'sh0086AE9F;
    weight_mem[ 154] = 32'shFFC08D97;
    weight_mem[ 155] = 32'shFEED1C52;
    weight_mem[ 156] = 32'shFE46CE80;
    weight_mem[ 157] = 32'sh02388EF0;
    weight_mem[ 158] = 32'shFBFF4EB0;
    weight_mem[ 159] = 32'sh0070B59D;
    weight_mem[ 160] = 32'shFAF4A780;
    weight_mem[ 161] = 32'shFDC9E1F8;
    weight_mem[ 162] = 32'shFCDDE3FC;
    weight_mem[ 163] = 32'sh01AD3B76;
    weight_mem[ 164] = 32'sh010AE908;
    weight_mem[ 165] = 32'sh01952CBC;
    weight_mem[ 166] = 32'shFC124BDC;
    weight_mem[ 167] = 32'sh091BA4E0;
    weight_mem[ 168] = 32'sh019212F2;
    weight_mem[ 169] = 32'sh00D8BE53;
    weight_mem[ 170] = 32'shFD4A60FC;
    weight_mem[ 171] = 32'sh00F1DB7A;
    weight_mem[ 172] = 32'sh03F7B388;
    weight_mem[ 173] = 32'shF85F0038;
    weight_mem[ 174] = 32'sh01EF8964;
    weight_mem[ 175] = 32'shFFAD902E;
    weight_mem[ 176] = 32'sh01F66E80;
    weight_mem[ 177] = 32'shFC1DADFC;
    weight_mem[ 178] = 32'shFD387970;
    weight_mem[ 179] = 32'shFE27C0B2;
    weight_mem[ 180] = 32'sh018CF15E;
    weight_mem[ 181] = 32'shFB9512D8;
    weight_mem[ 182] = 32'shFF147FB9;
    weight_mem[ 183] = 32'sh00203127;
    weight_mem[ 184] = 32'shF3CC97E0;
    weight_mem[ 185] = 32'sh0067D189;
    weight_mem[ 186] = 32'shFCB908C4;
    weight_mem[ 187] = 32'shFD58B968;
    weight_mem[ 188] = 32'shF49AE670;
    weight_mem[ 189] = 32'sh0A53ACE0;
    weight_mem[ 190] = 32'shFB199558;
    weight_mem[ 191] = 32'shFE2188D8;
    weight_mem[ 192] = 32'shFADD4768;
    weight_mem[ 193] = 32'shFB60FC50;
    weight_mem[ 194] = 32'sh0208A070;
    weight_mem[ 195] = 32'sh05130B60;
    weight_mem[ 196] = 32'shFD590ED4;
    weight_mem[ 197] = 32'shFF44B52A;
    weight_mem[ 198] = 32'sh02CDE06C;
    weight_mem[ 199] = 32'shFB00E660;
    weight_mem[ 200] = 32'shFC99BBC0;
    weight_mem[ 201] = 32'sh00E013BB;
    weight_mem[ 202] = 32'sh018BA08A;
    weight_mem[ 203] = 32'sh028AC924;
    weight_mem[ 204] = 32'sh009A0DDB;
    weight_mem[ 205] = 32'shFDE4C238;
    weight_mem[ 206] = 32'sh026EC620;
    weight_mem[ 207] = 32'shFD610078;
    weight_mem[ 208] = 32'sh052E4100;
    weight_mem[ 209] = 32'shFD3D6504;
    weight_mem[ 210] = 32'shFEB94AEE;
    weight_mem[ 211] = 32'shFE63235E;
    weight_mem[ 212] = 32'sh03B44170;
    weight_mem[ 213] = 32'shFCE3BD40;
    weight_mem[ 214] = 32'shFF9F01A4;
    weight_mem[ 215] = 32'sh014B534A;
    weight_mem[ 216] = 32'shFE8B1554;
    weight_mem[ 217] = 32'shFE4A467E;
    weight_mem[ 218] = 32'shFEEC60C0;
    weight_mem[ 219] = 32'shFA67DE88;
    weight_mem[ 220] = 32'shFDC8A24C;
    weight_mem[ 221] = 32'sh038CCFB4;
    weight_mem[ 222] = 32'shFFD344B6;
    weight_mem[ 223] = 32'sh029122AC;
    weight_mem[ 224] = 32'sh056240B8;
    weight_mem[ 225] = 32'sh001B15CB;
    weight_mem[ 226] = 32'shF966C370;
    weight_mem[ 227] = 32'sh04F78770;
    weight_mem[ 228] = 32'shFC2AFF48;
    weight_mem[ 229] = 32'sh0BD5F8C0;
    weight_mem[ 230] = 32'sh02279050;
    weight_mem[ 231] = 32'shFDF4CBE0;
    weight_mem[ 232] = 32'shFC64121C;
    weight_mem[ 233] = 32'sh0619BDC8;
    weight_mem[ 234] = 32'sh02453230;
    weight_mem[ 235] = 32'sh01A09E0A;
    weight_mem[ 236] = 32'sh0D3670F0;
    weight_mem[ 237] = 32'shFD5044F0;
    weight_mem[ 238] = 32'sh0267B924;
    weight_mem[ 239] = 32'sh03D7049C;
    weight_mem[ 240] = 32'shFE52EB58;
    weight_mem[ 241] = 32'sh00DD9B2F;
    weight_mem[ 242] = 32'sh06C9A0C0;
    weight_mem[ 243] = 32'shFC06036C;
    weight_mem[ 244] = 32'sh031A798C;
    weight_mem[ 245] = 32'sh007F36FE;
    weight_mem[ 246] = 32'sh01603AA8;
    weight_mem[ 247] = 32'shF1410DF0;
    weight_mem[ 248] = 32'shFB43AE78;
    weight_mem[ 249] = 32'shFCD9D6E4;
    weight_mem[ 250] = 32'sh029D77D4;
    weight_mem[ 251] = 32'sh02656F90;
    weight_mem[ 252] = 32'shFDFA3944;
    weight_mem[ 253] = 32'sh034259DC;
    weight_mem[ 254] = 32'sh0055D6AB;
    weight_mem[ 255] = 32'sh02C24564;
    weight_mem[ 256] = 32'sh00CA9350;
    weight_mem[ 257] = 32'sh00580E52;
    weight_mem[ 258] = 32'shFEDE7182;
    weight_mem[ 259] = 32'shFE25E218;
    weight_mem[ 260] = 32'shFFF81A78;
    weight_mem[ 261] = 32'sh019BDF1E;
    weight_mem[ 262] = 32'sh02209E28;
    weight_mem[ 263] = 32'sh013107F6;
    weight_mem[ 264] = 32'sh0144C578;
    weight_mem[ 265] = 32'shFABA6DF8;
    weight_mem[ 266] = 32'shFAF4D8C0;
    weight_mem[ 267] = 32'shFD9E8294;
    weight_mem[ 268] = 32'sh005FB5AA;
    weight_mem[ 269] = 32'shFC783C90;
    weight_mem[ 270] = 32'sh070D86B0;
    weight_mem[ 271] = 32'shFF7E7AE9;
    weight_mem[ 272] = 32'shFFE283D1;
    weight_mem[ 273] = 32'shFE4FB9F8;
    weight_mem[ 274] = 32'shFF60249C;
    weight_mem[ 275] = 32'shFD416234;
    weight_mem[ 276] = 32'shFEE43270;
    weight_mem[ 277] = 32'sh00450F3E;
    weight_mem[ 278] = 32'sh030BAE4C;
    weight_mem[ 279] = 32'shFE7C4D86;
    weight_mem[ 280] = 32'sh04335AF0;
    weight_mem[ 281] = 32'shFE6069CA;
    weight_mem[ 282] = 32'shFF1B54CE;
    weight_mem[ 283] = 32'sh02EF9630;
    weight_mem[ 284] = 32'shFFD8FB9A;
    weight_mem[ 285] = 32'shFB835090;
    weight_mem[ 286] = 32'shFF9A4E11;
    weight_mem[ 287] = 32'shFEF9F43A;
    weight_mem[ 288] = 32'sh04D505B0;
    weight_mem[ 289] = 32'shFFA646E6;
    weight_mem[ 290] = 32'sh00B0301A;
    weight_mem[ 291] = 32'sh02554264;
    weight_mem[ 292] = 32'sh022C6588;
    weight_mem[ 293] = 32'shFBDA6FC8;
    weight_mem[ 294] = 32'shFA2D1500;
    weight_mem[ 295] = 32'shFE87343E;
    weight_mem[ 296] = 32'sh02994C74;
    weight_mem[ 297] = 32'shFDB831DC;
    weight_mem[ 298] = 32'sh047C5F30;
    weight_mem[ 299] = 32'sh00AB53B5;
    weight_mem[ 300] = 32'sh00A597DD;
    weight_mem[ 301] = 32'shFE8EDCC4;
    weight_mem[ 302] = 32'sh04577890;
    weight_mem[ 303] = 32'shFE06217E;
    weight_mem[ 304] = 32'sh01F2000E;
    weight_mem[ 305] = 32'shFFDD551E;
    weight_mem[ 306] = 32'sh00A4EC6F;
    weight_mem[ 307] = 32'sh03011CC4;
    weight_mem[ 308] = 32'shFF79B606;
    weight_mem[ 309] = 32'shFF83F90F;
    weight_mem[ 310] = 32'shFD9F0B40;
    weight_mem[ 311] = 32'sh00AF9DF4;
    weight_mem[ 312] = 32'sh01933936;
    weight_mem[ 313] = 32'shFDE4C2D0;
    weight_mem[ 314] = 32'sh001CA384;
    weight_mem[ 315] = 32'shFEF935F4;
    weight_mem[ 316] = 32'sh0002C48F;
    weight_mem[ 317] = 32'sh00E361C5;
    weight_mem[ 318] = 32'shFCCCE3B0;
    weight_mem[ 319] = 32'shFFDC65DE;
    weight_mem[ 320] = 32'sh030931CC;
    weight_mem[ 321] = 32'shFEA92ADA;
    weight_mem[ 322] = 32'shFC6035AC;
    weight_mem[ 323] = 32'sh01945F16;
    weight_mem[ 324] = 32'sh01FCCCDE;
    weight_mem[ 325] = 32'sh026591F8;
    weight_mem[ 326] = 32'sh08A1E780;
    weight_mem[ 327] = 32'shF8B4E1B0;
    weight_mem[ 328] = 32'sh03F46928;
    weight_mem[ 329] = 32'shFFE13B44;
    weight_mem[ 330] = 32'sh040E0630;
    weight_mem[ 331] = 32'shFC290E00;
    weight_mem[ 332] = 32'sh03841F7C;
    weight_mem[ 333] = 32'shFF0CE712;
    weight_mem[ 334] = 32'sh04ED2A08;
    weight_mem[ 335] = 32'shFEBEAA98;
    weight_mem[ 336] = 32'shFC40F9E8;
    weight_mem[ 337] = 32'sh03690510;
    weight_mem[ 338] = 32'shFC8CD93C;
    weight_mem[ 339] = 32'shFF891EF7;
    weight_mem[ 340] = 32'sh057F82C0;
    weight_mem[ 341] = 32'sh02751C10;
    weight_mem[ 342] = 32'sh016A4492;
    weight_mem[ 343] = 32'sh00DDE65E;
    weight_mem[ 344] = 32'sh070789F8;
    weight_mem[ 345] = 32'shFC8C2EFC;
    weight_mem[ 346] = 32'sh00E67D51;
    weight_mem[ 347] = 32'sh034C11B8;
    weight_mem[ 348] = 32'shFB460E48;
    weight_mem[ 349] = 32'shFEE04828;
    weight_mem[ 350] = 32'sh01BC1A92;
    weight_mem[ 351] = 32'sh048E66E8;
    weight_mem[ 352] = 32'sh00C6D898;
    weight_mem[ 353] = 32'sh00112DFA;
    weight_mem[ 354] = 32'shFF325EAF;
    weight_mem[ 355] = 32'shFF3A3FE2;
    weight_mem[ 356] = 32'shFD63E480;
    weight_mem[ 357] = 32'sh0275ED58;
    weight_mem[ 358] = 32'sh03DF0DA4;
    weight_mem[ 359] = 32'sh024110D0;
    weight_mem[ 360] = 32'shFCD1673C;
    weight_mem[ 361] = 32'sh0372792C;
    weight_mem[ 362] = 32'shFA18F600;
    weight_mem[ 363] = 32'shFF927EEC;
    weight_mem[ 364] = 32'shFF302752;
    weight_mem[ 365] = 32'sh01670562;
    weight_mem[ 366] = 32'sh02BE6160;
    weight_mem[ 367] = 32'sh014D250A;
    weight_mem[ 368] = 32'shFF0D2A05;
    weight_mem[ 369] = 32'shFE2140A6;
    weight_mem[ 370] = 32'shFF27705F;
    weight_mem[ 371] = 32'shFDE659B4;
    weight_mem[ 372] = 32'sh00AC9CCE;
    weight_mem[ 373] = 32'shFDA553BC;
    weight_mem[ 374] = 32'sh01DF41E4;
    weight_mem[ 375] = 32'shFF49F1AE;
    weight_mem[ 376] = 32'shFB91FFB8;
    weight_mem[ 377] = 32'sh019475A2;
    weight_mem[ 378] = 32'shFF5C0956;
    weight_mem[ 379] = 32'shFEE415EE;
    weight_mem[ 380] = 32'sh011C071C;
    weight_mem[ 381] = 32'shFE682672;
    weight_mem[ 382] = 32'sh00BC6E26;
    weight_mem[ 383] = 32'shFFCC1B83;
    weight_mem[ 384] = 32'sh03A11C78;
    weight_mem[ 385] = 32'sh02C77078;
    weight_mem[ 386] = 32'sh013CDBC0;
    weight_mem[ 387] = 32'sh01067AA8;
    weight_mem[ 388] = 32'shF81E4DC0;
    weight_mem[ 389] = 32'shFE9F02B8;
    weight_mem[ 390] = 32'shFE6AE900;
    weight_mem[ 391] = 32'shFF83B4BA;
    weight_mem[ 392] = 32'shEFF041C0;
    weight_mem[ 393] = 32'shFE95503C;
    weight_mem[ 394] = 32'shFF1BF97C;
    weight_mem[ 395] = 32'shFE9D3EDE;
    weight_mem[ 396] = 32'sh011E89A0;
    weight_mem[ 397] = 32'sh03DE65D0;
    weight_mem[ 398] = 32'shFFFCD003;
    weight_mem[ 399] = 32'shFE163794;
    weight_mem[ 400] = 32'sh060613B8;
    weight_mem[ 401] = 32'sh01495D2A;
    weight_mem[ 402] = 32'shFD74BC68;
    weight_mem[ 403] = 32'sh000DF40B;
    weight_mem[ 404] = 32'shF8FD6870;
    weight_mem[ 405] = 32'sh05A39510;
    weight_mem[ 406] = 32'shFE0DC2BC;
    weight_mem[ 407] = 32'shFFCC2419;
    weight_mem[ 408] = 32'sh062EC5E8;
    weight_mem[ 409] = 32'shFD9FE074;
    weight_mem[ 410] = 32'sh03D89290;
    weight_mem[ 411] = 32'shFF475AC9;
    weight_mem[ 412] = 32'sh013AD5E4;
    weight_mem[ 413] = 32'shFD0F4348;
    weight_mem[ 414] = 32'sh06A4A988;
    weight_mem[ 415] = 32'shFF109CF0;
    weight_mem[ 416] = 32'shFEDBE3A6;
    weight_mem[ 417] = 32'sh075E9DA8;
    weight_mem[ 418] = 32'sh05C919A0;
    weight_mem[ 419] = 32'sh00497430;
    weight_mem[ 420] = 32'shFDC950D0;
    weight_mem[ 421] = 32'shF4A36CB0;
    weight_mem[ 422] = 32'shFA1E3860;
    weight_mem[ 423] = 32'sh019B98A8;
    weight_mem[ 424] = 32'sh026283D4;
    weight_mem[ 425] = 32'sh008D8242;
    weight_mem[ 426] = 32'sh01468EE0;
    weight_mem[ 427] = 32'sh048F1838;
    weight_mem[ 428] = 32'shF8042F10;
    weight_mem[ 429] = 32'sh0F60EF10;
    weight_mem[ 430] = 32'shFCC4E1D0;
    weight_mem[ 431] = 32'shF82CA670;
    weight_mem[ 432] = 32'shFF883AEC;
    weight_mem[ 433] = 32'sh021B477C;
    weight_mem[ 434] = 32'sh08036150;
    weight_mem[ 435] = 32'sh0156B9A0;
    weight_mem[ 436] = 32'sh0395D068;
    weight_mem[ 437] = 32'shFC18E948;
    weight_mem[ 438] = 32'shFE6EDF28;
    weight_mem[ 439] = 32'shFB713390;
    weight_mem[ 440] = 32'sh055C7440;
    weight_mem[ 441] = 32'shFDBC82A8;
    weight_mem[ 442] = 32'shFED1AA70;
    weight_mem[ 443] = 32'sh02784724;
    weight_mem[ 444] = 32'sh0A8792F0;
    weight_mem[ 445] = 32'shF55D2280;
    weight_mem[ 446] = 32'shFDAD0FB8;
    weight_mem[ 447] = 32'sh04B6EB50;
    weight_mem[ 448] = 32'shF6A20050;
    weight_mem[ 449] = 32'sh00B30BCD;
    weight_mem[ 450] = 32'sh011A987E;
    weight_mem[ 451] = 32'sh00A29FD1;
    weight_mem[ 452] = 32'sh067AF1E0;
    weight_mem[ 453] = 32'shFDA00068;
    weight_mem[ 454] = 32'sh05D50C38;
    weight_mem[ 455] = 32'sh0409B388;
    weight_mem[ 456] = 32'shFD448558;
    weight_mem[ 457] = 32'shF622E1A0;
    weight_mem[ 458] = 32'sh09465140;
    weight_mem[ 459] = 32'shF772BE90;
    weight_mem[ 460] = 32'shFDC8B6D4;
    weight_mem[ 461] = 32'shF0091C90;
    weight_mem[ 462] = 32'shFF422FFD;
    weight_mem[ 463] = 32'sh02ABEE08;
    weight_mem[ 464] = 32'sh09B0BB90;
    weight_mem[ 465] = 32'shFF8EFB3D;
    weight_mem[ 466] = 32'shF9CD1550;
    weight_mem[ 467] = 32'sh045BC0F0;
    weight_mem[ 468] = 32'shFC545F70;
    weight_mem[ 469] = 32'sh01F194E4;
    weight_mem[ 470] = 32'shFFCC4C37;
    weight_mem[ 471] = 32'sh081269B0;
    weight_mem[ 472] = 32'shF3CEA3A0;
    weight_mem[ 473] = 32'shF719D4A0;
    weight_mem[ 474] = 32'sh068BABD8;
    weight_mem[ 475] = 32'shFEE4E96A;
    weight_mem[ 476] = 32'shF94D3478;
    weight_mem[ 477] = 32'sh0EFEC130;
    weight_mem[ 478] = 32'shED927740;
    weight_mem[ 479] = 32'shFAF9A4E8;
    weight_mem[ 480] = 32'sh032A5D30;
    weight_mem[ 481] = 32'sh009E3138;
    weight_mem[ 482] = 32'shFB576200;
    weight_mem[ 483] = 32'sh0563AF90;
    weight_mem[ 484] = 32'sh01F268E4;
    weight_mem[ 485] = 32'sh09CA5290;
    weight_mem[ 486] = 32'sh00B7EB47;
    weight_mem[ 487] = 32'shFFC13A24;
    weight_mem[ 488] = 32'sh05121248;
    weight_mem[ 489] = 32'shFA1DA728;
    weight_mem[ 490] = 32'sh03131490;
    weight_mem[ 491] = 32'sh03B6043C;
    weight_mem[ 492] = 32'sh01FC2684;
    weight_mem[ 493] = 32'sh0132167C;
    weight_mem[ 494] = 32'sh01A29128;
    weight_mem[ 495] = 32'sh00DB5AF8;
    weight_mem[ 496] = 32'shFE1AD45E;
    weight_mem[ 497] = 32'sh0183CA30;
    weight_mem[ 498] = 32'shFF313069;
    weight_mem[ 499] = 32'shFB3D3E90;
    weight_mem[ 500] = 32'sh01E91D12;
    weight_mem[ 501] = 32'shFD64E638;
    weight_mem[ 502] = 32'shFFE28720;
    weight_mem[ 503] = 32'sh008EA628;
    weight_mem[ 504] = 32'sh04AE70F8;
    weight_mem[ 505] = 32'shFBFAEEF8;
    weight_mem[ 506] = 32'shFC0054A4;
    weight_mem[ 507] = 32'sh007C9FDB;
    weight_mem[ 508] = 32'sh02D28804;
    weight_mem[ 509] = 32'shFDF8F87C;
    weight_mem[ 510] = 32'shF90F5468;
    weight_mem[ 511] = 32'shFFD187BE;
    weight_mem[ 512] = 32'sh01C59CBE;
    weight_mem[ 513] = 32'shFF726FB9;
    weight_mem[ 514] = 32'shFB862340;
    weight_mem[ 515] = 32'shFD79B334;
    weight_mem[ 516] = 32'shFEDF82EA;
    weight_mem[ 517] = 32'sh02089E84;
    weight_mem[ 518] = 32'shFF7B9E0D;
    weight_mem[ 519] = 32'sh0265D8F8;
    weight_mem[ 520] = 32'sh01E7F838;
    weight_mem[ 521] = 32'sh0067FBCF;
    weight_mem[ 522] = 32'shF8887A90;
    weight_mem[ 523] = 32'shFFFB7EF3;
    weight_mem[ 524] = 32'shFFFA6545;
    weight_mem[ 525] = 32'sh03CD1B20;
    weight_mem[ 526] = 32'sh04E2ADC0;
    weight_mem[ 527] = 32'shFFE5BEEF;
    weight_mem[ 528] = 32'sh006B6DDC;
    weight_mem[ 529] = 32'sh021FEF94;
    weight_mem[ 530] = 32'sh034D7600;
    weight_mem[ 531] = 32'shFE5B21C6;
    weight_mem[ 532] = 32'shFD62B914;
    weight_mem[ 533] = 32'sh007A1364;
    weight_mem[ 534] = 32'sh0216C32C;
    weight_mem[ 535] = 32'shFDDE4E1C;
    weight_mem[ 536] = 32'shFFF802B0;
    weight_mem[ 537] = 32'sh036B4EF0;
    weight_mem[ 538] = 32'shFE7A5246;
    weight_mem[ 539] = 32'sh0199F44E;
    weight_mem[ 540] = 32'shFF0C209F;
    weight_mem[ 541] = 32'shFF7FC24A;
    weight_mem[ 542] = 32'sh00FB2B3A;
    weight_mem[ 543] = 32'shFFCBDB64;
    weight_mem[ 544] = 32'shFDDA7A58;
    weight_mem[ 545] = 32'sh02918530;
    weight_mem[ 546] = 32'shFE8D931C;
    weight_mem[ 547] = 32'shFB478BD0;
    weight_mem[ 548] = 32'shFFB5AE26;
    weight_mem[ 549] = 32'shFF3B69A0;
    weight_mem[ 550] = 32'shF20918B0;
    weight_mem[ 551] = 32'sh032690BC;
    weight_mem[ 552] = 32'shFD696784;
    weight_mem[ 553] = 32'shFA606988;
    weight_mem[ 554] = 32'shFF29AE4E;
    weight_mem[ 555] = 32'shFFB4DDCE;
    weight_mem[ 556] = 32'shFFCCB98C;
    weight_mem[ 557] = 32'shFFDC46B0;
    weight_mem[ 558] = 32'shFEBBC63C;
    weight_mem[ 559] = 32'sh016F9214;
    weight_mem[ 560] = 32'sh00293826;
    weight_mem[ 561] = 32'shFF1BD1C9;
    weight_mem[ 562] = 32'sh01E0952C;
    weight_mem[ 563] = 32'sh017277A6;
    weight_mem[ 564] = 32'shFEAD58BE;
    weight_mem[ 565] = 32'sh001112DF;
    weight_mem[ 566] = 32'shF9B405F0;
    weight_mem[ 567] = 32'shFC5AB110;
    weight_mem[ 568] = 32'shFEB5802A;
    weight_mem[ 569] = 32'shFC8B7CB4;
    weight_mem[ 570] = 32'sh0488B1D8;
    weight_mem[ 571] = 32'sh0248442C;
    weight_mem[ 572] = 32'sh05775760;
    weight_mem[ 573] = 32'shFADF1798;
    weight_mem[ 574] = 32'shFAA29B78;
    weight_mem[ 575] = 32'shFF2D7532;
    weight_mem[ 576] = 32'shFF1BEA2B;
    weight_mem[ 577] = 32'sh06F686F0;
    weight_mem[ 578] = 32'sh07F3B9F0;
    weight_mem[ 579] = 32'sh018E11B0;
    weight_mem[ 580] = 32'shFE39864C;
    weight_mem[ 581] = 32'shFD1BB810;
    weight_mem[ 582] = 32'shFB3094C0;
    weight_mem[ 583] = 32'shFE868736;
    weight_mem[ 584] = 32'sh02CE62D0;
    weight_mem[ 585] = 32'sh00699BC0;
    weight_mem[ 586] = 32'sh0489A820;
    weight_mem[ 587] = 32'sh03A0B340;
    weight_mem[ 588] = 32'shF5AAFE20;
    weight_mem[ 589] = 32'sh0EEF5600;
    weight_mem[ 590] = 32'shFA0F2E38;
    weight_mem[ 591] = 32'shF8A2A350;
    weight_mem[ 592] = 32'shFF1A9AEE;
    weight_mem[ 593] = 32'sh0591C7C8;
    weight_mem[ 594] = 32'sh05EBA8A0;
    weight_mem[ 595] = 32'shF8227078;
    weight_mem[ 596] = 32'sh0480B948;
    weight_mem[ 597] = 32'shFB9C0D98;
    weight_mem[ 598] = 32'sh0111249A;
    weight_mem[ 599] = 32'shFE66F8E2;
    weight_mem[ 600] = 32'sh07932320;
    weight_mem[ 601] = 32'shFDA7E9C8;
    weight_mem[ 602] = 32'shFDF70E44;
    weight_mem[ 603] = 32'sh00DD1FF5;
    weight_mem[ 604] = 32'sh090A2410;
    weight_mem[ 605] = 32'shF65124E0;
    weight_mem[ 606] = 32'sh0085E770;
    weight_mem[ 607] = 32'sh04F3A908;
    weight_mem[ 608] = 32'sh035BBD14;
    weight_mem[ 609] = 32'sh04926018;
    weight_mem[ 610] = 32'shFF3B3096;
    weight_mem[ 611] = 32'shFFBC5717;
    weight_mem[ 612] = 32'sh00E30275;
    weight_mem[ 613] = 32'shFD633D90;
    weight_mem[ 614] = 32'shFFB53A8A;
    weight_mem[ 615] = 32'shFDE2A014;
    weight_mem[ 616] = 32'shFF47AF41;
    weight_mem[ 617] = 32'shFF9B84FC;
    weight_mem[ 618] = 32'sh04E76798;
    weight_mem[ 619] = 32'sh0002F64A;
    weight_mem[ 620] = 32'shFF83458C;
    weight_mem[ 621] = 32'sh00598DB9;
    weight_mem[ 622] = 32'sh063AD1E0;
    weight_mem[ 623] = 32'shFEA00710;
    weight_mem[ 624] = 32'sh0203F5E8;
    weight_mem[ 625] = 32'sh04CE3488;
    weight_mem[ 626] = 32'sh067F14D8;
    weight_mem[ 627] = 32'sh0119804A;
    weight_mem[ 628] = 32'shFD2F6814;
    weight_mem[ 629] = 32'sh06B5E2E8;
    weight_mem[ 630] = 32'shFE650B1A;
    weight_mem[ 631] = 32'shFD023DFC;
    weight_mem[ 632] = 32'shFB422E80;
    weight_mem[ 633] = 32'shF9E566E0;
    weight_mem[ 634] = 32'sh066FF670;
    weight_mem[ 635] = 32'sh013D9A38;
    weight_mem[ 636] = 32'sh04F5A7D0;
    weight_mem[ 637] = 32'sh0082631A;
    weight_mem[ 638] = 32'shF60EEAD0;
    weight_mem[ 639] = 32'sh0056C6B2;
    weight_mem[ 640] = 32'shFD24AE20;
    weight_mem[ 641] = 32'shFCCB5914;
    weight_mem[ 642] = 32'sh0259FE50;
    weight_mem[ 643] = 32'shFED139FA;
    weight_mem[ 644] = 32'sh02B4548C;
    weight_mem[ 645] = 32'shF97A8708;
    weight_mem[ 646] = 32'shFFFB0C6A;
    weight_mem[ 647] = 32'sh037621B8;
    weight_mem[ 648] = 32'shFD8FEF48;
    weight_mem[ 649] = 32'sh024CE8D0;
    weight_mem[ 650] = 32'sh00F8F893;
    weight_mem[ 651] = 32'shFDC83294;
    weight_mem[ 652] = 32'sh00D544B0;
    weight_mem[ 653] = 32'shFF8CB2E0;
    weight_mem[ 654] = 32'shFBB5ED70;
    weight_mem[ 655] = 32'sh00838BB6;
    weight_mem[ 656] = 32'sh0543B910;
    weight_mem[ 657] = 32'sh03611748;
    weight_mem[ 658] = 32'sh041A6120;
    weight_mem[ 659] = 32'sh049F99D8;
    weight_mem[ 660] = 32'shF80239B0;
    weight_mem[ 661] = 32'shFCBC6F0C;
    weight_mem[ 662] = 32'shFC7C480C;
    weight_mem[ 663] = 32'shFE439B8E;
    weight_mem[ 664] = 32'shFB3B1728;
    weight_mem[ 665] = 32'sh009B711F;
    weight_mem[ 666] = 32'shFDF316D0;
    weight_mem[ 667] = 32'shFAEB9118;
    weight_mem[ 668] = 32'sh0B302DD0;
    weight_mem[ 669] = 32'sh00617556;
    weight_mem[ 670] = 32'shFA3AA898;
    weight_mem[ 671] = 32'shFFE3BA44;
    weight_mem[ 672] = 32'shFD1AB42C;
    weight_mem[ 673] = 32'sh00691D33;
    weight_mem[ 674] = 32'shFE6D7E4C;
    weight_mem[ 675] = 32'sh0AC7D8C0;
    weight_mem[ 676] = 32'shFE4C7896;
    weight_mem[ 677] = 32'sh046FF540;
    weight_mem[ 678] = 32'shFC0C5D28;
    weight_mem[ 679] = 32'sh0237A4D8;
    weight_mem[ 680] = 32'shFA7B0298;
    weight_mem[ 681] = 32'shFB6D7730;
    weight_mem[ 682] = 32'sh0445DE10;
    weight_mem[ 683] = 32'sh009C4951;
    weight_mem[ 684] = 32'sh012A5762;
    weight_mem[ 685] = 32'sh009C5DD9;
    weight_mem[ 686] = 32'sh00D21F4C;
    weight_mem[ 687] = 32'sh00E4FC57;
    weight_mem[ 688] = 32'sh042A0FE8;
    weight_mem[ 689] = 32'shF8B72740;
    weight_mem[ 690] = 32'sh029A0D5C;
    weight_mem[ 691] = 32'shFBA4C7A8;
    weight_mem[ 692] = 32'sh00CB2FDE;
    weight_mem[ 693] = 32'shF69A1040;
    weight_mem[ 694] = 32'shFC545500;
    weight_mem[ 695] = 32'shFDB0725C;
    weight_mem[ 696] = 32'sh01CDE144;
    weight_mem[ 697] = 32'shFBA09470;
    weight_mem[ 698] = 32'shFE05D286;
    weight_mem[ 699] = 32'shFA4A6548;
    weight_mem[ 700] = 32'shFBA6B1A0;
    weight_mem[ 701] = 32'shFDAA3C4C;
    weight_mem[ 702] = 32'shFC513668;
    weight_mem[ 703] = 32'shFFAE1170;
    weight_mem[ 704] = 32'sh04E20CE8;
    weight_mem[ 705] = 32'shFD9920A4;
    weight_mem[ 706] = 32'shFFB6AAAD;
    weight_mem[ 707] = 32'shFDD057D0;
    weight_mem[ 708] = 32'shFB26CDE0;
    weight_mem[ 709] = 32'sh04B6D748;
    weight_mem[ 710] = 32'shFC7D46A4;
    weight_mem[ 711] = 32'shFD30C654;
    weight_mem[ 712] = 32'sh01D9519E;
    weight_mem[ 713] = 32'shFE923CA8;
    weight_mem[ 714] = 32'sh0082B4A7;
    weight_mem[ 715] = 32'sh026248A0;
    weight_mem[ 716] = 32'sh020DAEB4;
    weight_mem[ 717] = 32'sh05BEBA80;
    weight_mem[ 718] = 32'shFC7B43B4;
    weight_mem[ 719] = 32'sh025F6078;
    weight_mem[ 720] = 32'shFC0C5848;
    weight_mem[ 721] = 32'sh04E16F68;
    weight_mem[ 722] = 32'sh00FFB099;
    weight_mem[ 723] = 32'shFA9ADF20;
    weight_mem[ 724] = 32'shFE35CD2C;
    weight_mem[ 725] = 32'sh054A11A8;
    weight_mem[ 726] = 32'shFE8FB91C;
    weight_mem[ 727] = 32'shFF231B98;
    weight_mem[ 728] = 32'sh062BC270;
    weight_mem[ 729] = 32'sh026E952C;
    weight_mem[ 730] = 32'shFF2BF491;
    weight_mem[ 731] = 32'sh060B7EA0;
    weight_mem[ 732] = 32'sh04844C08;
    weight_mem[ 733] = 32'shFF4162FD;
    weight_mem[ 734] = 32'sh02853A4C;
    weight_mem[ 735] = 32'shFE68CAEE;
    weight_mem[ 736] = 32'sh051D3A90;
    weight_mem[ 737] = 32'sh003C34B6;
    weight_mem[ 738] = 32'shFF915F58;
    weight_mem[ 739] = 32'sh0083895B;
    weight_mem[ 740] = 32'sh0375DF54;
    weight_mem[ 741] = 32'shFAB77D68;
    weight_mem[ 742] = 32'shF7FA1BD0;
    weight_mem[ 743] = 32'sh016B7432;
    weight_mem[ 744] = 32'sh04790B68;
    weight_mem[ 745] = 32'shFADD1130;
    weight_mem[ 746] = 32'sh04554F60;
    weight_mem[ 747] = 32'sh006EF71F;
    weight_mem[ 748] = 32'shFA12BDD8;
    weight_mem[ 749] = 32'sh029757A8;
    weight_mem[ 750] = 32'sh0379145C;
    weight_mem[ 751] = 32'sh03C4552C;
    weight_mem[ 752] = 32'shFCC6797C;
    weight_mem[ 753] = 32'sh087496D0;
    weight_mem[ 754] = 32'shFFCFA2FE;
    weight_mem[ 755] = 32'sh0163EDD2;
    weight_mem[ 756] = 32'shFAEB16F0;
    weight_mem[ 757] = 32'shFE037CAE;
    weight_mem[ 758] = 32'shFEED86CA;
    weight_mem[ 759] = 32'sh07F929C8;
    weight_mem[ 760] = 32'sh0399EFE8;
    weight_mem[ 761] = 32'sh01A347AC;
    weight_mem[ 762] = 32'sh02670734;
    weight_mem[ 763] = 32'shFB9B1D20;
    weight_mem[ 764] = 32'sh00F64C40;
    weight_mem[ 765] = 32'shFDD557D4;
    weight_mem[ 766] = 32'shFE15AADC;
    weight_mem[ 767] = 32'sh023D24C8;
    weight_mem[ 768] = 32'sh008B78B1;
    weight_mem[ 769] = 32'sh00B465B6;
    weight_mem[ 770] = 32'sh03CE3328;
    weight_mem[ 771] = 32'shFA1C6F78;
    weight_mem[ 772] = 32'sh04D35408;
    weight_mem[ 773] = 32'shFC664DA4;
    weight_mem[ 774] = 32'sh01DD810C;
    weight_mem[ 775] = 32'sh02C26A34;
    weight_mem[ 776] = 32'sh03DE697C;
    weight_mem[ 777] = 32'sh035A589C;
    weight_mem[ 778] = 32'shFDFE60FC;
    weight_mem[ 779] = 32'shFDC5A014;
    weight_mem[ 780] = 32'shFF0310D0;
    weight_mem[ 781] = 32'sh0147421E;
    weight_mem[ 782] = 32'sh057EDE40;
    weight_mem[ 783] = 32'shFCE90644;
    weight_mem[ 784] = 32'sh00C1E375;
    weight_mem[ 785] = 32'shFE4BA3BA;
    weight_mem[ 786] = 32'sh02AA5274;
    weight_mem[ 787] = 32'sh005BC7E4;
    weight_mem[ 788] = 32'shFE8D2B02;
    weight_mem[ 789] = 32'shFDBCE028;
    weight_mem[ 790] = 32'shFB08A4D8;
    weight_mem[ 791] = 32'shFF9CD922;
    weight_mem[ 792] = 32'shF90EC460;
    weight_mem[ 793] = 32'shFF3EFFFD;
    weight_mem[ 794] = 32'shFE304C6C;
    weight_mem[ 795] = 32'sh0022E85C;
    weight_mem[ 796] = 32'sh04E8C4F8;
    weight_mem[ 797] = 32'sh0057F81A;
    weight_mem[ 798] = 32'shFC44646C;
    weight_mem[ 799] = 32'sh02ACF778;
    weight_mem[ 800] = 32'shFFC823F1;
    weight_mem[ 801] = 32'sh01BE9600;
    weight_mem[ 802] = 32'shFE4D7B5E;
    weight_mem[ 803] = 32'sh077E77E0;
    weight_mem[ 804] = 32'shFF25D5F9;
    weight_mem[ 805] = 32'shFC17B1E8;
    weight_mem[ 806] = 32'sh024CA30C;
    weight_mem[ 807] = 32'shFE307972;
    weight_mem[ 808] = 32'shFF19369D;
    weight_mem[ 809] = 32'sh01C94C8A;
    weight_mem[ 810] = 32'sh00D7B749;
    weight_mem[ 811] = 32'sh03028618;
    weight_mem[ 812] = 32'shFE865EB6;
    weight_mem[ 813] = 32'sh01357B1E;
    weight_mem[ 814] = 32'sh01069B8A;
    weight_mem[ 815] = 32'shFDCA41E8;
    weight_mem[ 816] = 32'shFF2E57C1;
    weight_mem[ 817] = 32'sh005B73DD;
    weight_mem[ 818] = 32'shFD0E80D4;
    weight_mem[ 819] = 32'sh04D30768;
    weight_mem[ 820] = 32'shFAB25348;
    weight_mem[ 821] = 32'shFE1DD066;
    weight_mem[ 822] = 32'sh0215B2D4;
    weight_mem[ 823] = 32'sh043718A8;
    weight_mem[ 824] = 32'sh003BACE5;
    weight_mem[ 825] = 32'shFD88F2C4;
    weight_mem[ 826] = 32'shF998BED0;
    weight_mem[ 827] = 32'shF7169B30;
    weight_mem[ 828] = 32'shFDFCB60C;
    weight_mem[ 829] = 32'sh015DF96C;
    weight_mem[ 830] = 32'sh027A335C;
    weight_mem[ 831] = 32'sh027D44E8;
    weight_mem[ 832] = 32'shFE9CD9A2;
    weight_mem[ 833] = 32'shFE33B7A0;
    weight_mem[ 834] = 32'sh0130FB7C;
    weight_mem[ 835] = 32'shFD3FCCDC;
    weight_mem[ 836] = 32'sh06704478;
    weight_mem[ 837] = 32'shFCFCF8F4;
    weight_mem[ 838] = 32'shFCAC7798;
    weight_mem[ 839] = 32'sh04CC0000;
    weight_mem[ 840] = 32'sh05C486C8;
    weight_mem[ 841] = 32'shF84F0D70;
    weight_mem[ 842] = 32'sh021A7BD0;
    weight_mem[ 843] = 32'sh00B33DB8;
    weight_mem[ 844] = 32'shFABE4B68;
    weight_mem[ 845] = 32'sh00007AFC;
    weight_mem[ 846] = 32'sh045CFE60;
    weight_mem[ 847] = 32'sh04A10B30;
    weight_mem[ 848] = 32'sh01A56ECC;
    weight_mem[ 849] = 32'sh02B6BAE8;
    weight_mem[ 850] = 32'sh09387300;
    weight_mem[ 851] = 32'sh013CAB66;
    weight_mem[ 852] = 32'sh02C9885C;
    weight_mem[ 853] = 32'shFD714EB0;
    weight_mem[ 854] = 32'sh01F2F0A4;
    weight_mem[ 855] = 32'shFE017A54;
    weight_mem[ 856] = 32'sh08C5D9F0;
    weight_mem[ 857] = 32'shFE059B5A;
    weight_mem[ 858] = 32'shFCE29E38;
    weight_mem[ 859] = 32'shFE654698;
    weight_mem[ 860] = 32'shFE550FD2;
    weight_mem[ 861] = 32'shFEB150B0;
    weight_mem[ 862] = 32'sh008566CF;
    weight_mem[ 863] = 32'shFED531A8;
    weight_mem[ 864] = 32'sh0C0C1CD0;
    weight_mem[ 865] = 32'shFE93602C;
    weight_mem[ 866] = 32'shFF20AFC5;
    weight_mem[ 867] = 32'shFCCA2814;
    weight_mem[ 868] = 32'shF7B1E330;
    weight_mem[ 869] = 32'sh00B56419;
    weight_mem[ 870] = 32'shF906CA80;
    weight_mem[ 871] = 32'shFD506134;
    weight_mem[ 872] = 32'shFFB375AA;
    weight_mem[ 873] = 32'sh041DCB70;
    weight_mem[ 874] = 32'shF6838920;
    weight_mem[ 875] = 32'sh08BD1DB0;
    weight_mem[ 876] = 32'sh02E958BC;
    weight_mem[ 877] = 32'sh0F427650;
    weight_mem[ 878] = 32'shFC94E03C;
    weight_mem[ 879] = 32'shFD6EC730;
    weight_mem[ 880] = 32'shF6DD63F0;
    weight_mem[ 881] = 32'shFC6F40D0;
    weight_mem[ 882] = 32'sh066C9EF0;
    weight_mem[ 883] = 32'shFD09E9A8;
    weight_mem[ 884] = 32'sh043CF818;
    weight_mem[ 885] = 32'shFEFBB40E;
    weight_mem[ 886] = 32'shFDE2EFA4;
    weight_mem[ 887] = 32'shF79CC3D0;
    weight_mem[ 888] = 32'sh0EFD9360;
    weight_mem[ 889] = 32'sh0B5477F0;
    weight_mem[ 890] = 32'shF9B1A498;
    weight_mem[ 891] = 32'sh020AA3A0;
    weight_mem[ 892] = 32'sh142A6F60;
    weight_mem[ 893] = 32'shF0C5E780;
    weight_mem[ 894] = 32'sh08655BE0;
    weight_mem[ 895] = 32'sh04F92648;
    weight_mem[ 896] = 32'shFA098330;
    weight_mem[ 897] = 32'sh00EC74C4;
    weight_mem[ 898] = 32'sh00B0EDA6;
    weight_mem[ 899] = 32'sh0546D6F8;
    weight_mem[ 900] = 32'sh01026A58;
    weight_mem[ 901] = 32'shFFE7EBF6;
    weight_mem[ 902] = 32'sh01213D0E;
    weight_mem[ 903] = 32'shFCE1FD14;
    weight_mem[ 904] = 32'shFFAFF2C8;
    weight_mem[ 905] = 32'shFCD69C50;
    weight_mem[ 906] = 32'sh03E6F638;
    weight_mem[ 907] = 32'shFDAA2980;
    weight_mem[ 908] = 32'shFDB891F8;
    weight_mem[ 909] = 32'sh04F359D0;
    weight_mem[ 910] = 32'shF9C56F90;
    weight_mem[ 911] = 32'sh01BD4D12;
    weight_mem[ 912] = 32'shFE11200A;
    weight_mem[ 913] = 32'sh0140E300;
    weight_mem[ 914] = 32'sh0A674580;
    weight_mem[ 915] = 32'shFE6AB9F4;
    weight_mem[ 916] = 32'shFD9C3E2C;
    weight_mem[ 917] = 32'shFEC018F0;
    weight_mem[ 918] = 32'sh0007AF56;
    weight_mem[ 919] = 32'sh00338001;
    weight_mem[ 920] = 32'sh0059D82A;
    weight_mem[ 921] = 32'shFF82C0A1;
    weight_mem[ 922] = 32'shFF08CA29;
    weight_mem[ 923] = 32'shFADEDFB8;
    weight_mem[ 924] = 32'shFE0ED04E;
    weight_mem[ 925] = 32'shFE682FEE;
    weight_mem[ 926] = 32'shFFC2CBEF;
    weight_mem[ 927] = 32'sh03810CEC;
    weight_mem[ 928] = 32'sh05F5E4D0;
    weight_mem[ 929] = 32'sh016A0B48;
    weight_mem[ 930] = 32'shFDC411D4;
    weight_mem[ 931] = 32'sh034B9B9C;
    weight_mem[ 932] = 32'shF920A638;
    weight_mem[ 933] = 32'shFE14267C;
    weight_mem[ 934] = 32'sh011DB348;
    weight_mem[ 935] = 32'shFE076044;
    weight_mem[ 936] = 32'shFF7402AD;
    weight_mem[ 937] = 32'shFF5FE237;
    weight_mem[ 938] = 32'sh040BDC58;
    weight_mem[ 939] = 32'sh018A9C02;
    weight_mem[ 940] = 32'sh04A13A38;
    weight_mem[ 941] = 32'shFF3DE3F3;
    weight_mem[ 942] = 32'shF73931C0;
    weight_mem[ 943] = 32'sh00FEBB7F;
    weight_mem[ 944] = 32'shF7388740;
    weight_mem[ 945] = 32'shFBABFF98;
    weight_mem[ 946] = 32'shFE33342A;
    weight_mem[ 947] = 32'sh04647E18;
    weight_mem[ 948] = 32'sh048718D8;
    weight_mem[ 949] = 32'shFD6B05A8;
    weight_mem[ 950] = 32'sh01D50012;
    weight_mem[ 951] = 32'shFB9CE508;
    weight_mem[ 952] = 32'sh02DFB2D4;
    weight_mem[ 953] = 32'sh048CF2B8;
    weight_mem[ 954] = 32'sh028791BC;
    weight_mem[ 955] = 32'sh00D1199C;
    weight_mem[ 956] = 32'sh00F73BA8;
    weight_mem[ 957] = 32'shFFE48870;
    weight_mem[ 958] = 32'sh0579D530;
    weight_mem[ 959] = 32'sh037F2AB0;
    weight_mem[ 960] = 32'shFEE712DA;
    weight_mem[ 961] = 32'sh077EBC60;
    weight_mem[ 962] = 32'sh03105580;
    weight_mem[ 963] = 32'sh0124E23E;
    weight_mem[ 964] = 32'shFF06C1D9;
    weight_mem[ 965] = 32'sh05634788;
    weight_mem[ 966] = 32'sh054D0700;
    weight_mem[ 967] = 32'sh02C5CD08;
    weight_mem[ 968] = 32'sh0228B6B0;
    weight_mem[ 969] = 32'shFD35B1F0;
    weight_mem[ 970] = 32'shFFCA3698;
    weight_mem[ 971] = 32'shFD1C0094;
    weight_mem[ 972] = 32'shF81AAC98;
    weight_mem[ 973] = 32'sh06184BD8;
    weight_mem[ 974] = 32'sh06D43B80;
    weight_mem[ 975] = 32'shF7198480;
    weight_mem[ 976] = 32'shFF897358;
    weight_mem[ 977] = 32'sh028BB814;
    weight_mem[ 978] = 32'sh00158199;
    weight_mem[ 979] = 32'shF8315208;
    weight_mem[ 980] = 32'sh00FDABD1;
    weight_mem[ 981] = 32'shF9E454B0;
    weight_mem[ 982] = 32'shFC56B138;
    weight_mem[ 983] = 32'sh0855D090;
    weight_mem[ 984] = 32'sh00FC5892;
    weight_mem[ 985] = 32'shFCE1D730;
    weight_mem[ 986] = 32'shFE39B95E;
    weight_mem[ 987] = 32'sh007ED6C6;
    weight_mem[ 988] = 32'sh02D98860;
    weight_mem[ 989] = 32'shFC316994;
    weight_mem[ 990] = 32'shFA574AF8;
    weight_mem[ 991] = 32'sh05ED3CF8;
    weight_mem[ 992] = 32'shFB586A30;
    weight_mem[ 993] = 32'sh013E8BF0;
    weight_mem[ 994] = 32'shFE3EE9D2;
    weight_mem[ 995] = 32'sh021A0D1C;
    weight_mem[ 996] = 32'shFF11E930;
    weight_mem[ 997] = 32'sh00F5E7CD;
    weight_mem[ 998] = 32'sh00EC2C22;
    weight_mem[ 999] = 32'shFDD7BE68;
    weight_mem[1000] = 32'shFEEEB70E;
    weight_mem[1001] = 32'sh037008C0;
    weight_mem[1002] = 32'shFBE07A60;
    weight_mem[1003] = 32'shFFA15364;
    weight_mem[1004] = 32'sh00FDCEFE;
    weight_mem[1005] = 32'sh0277ACEC;
    weight_mem[1006] = 32'shFF7062AA;
    weight_mem[1007] = 32'shFF83B7F6;
    weight_mem[1008] = 32'shFF21ACC8;
    weight_mem[1009] = 32'sh0143EFE0;
    weight_mem[1010] = 32'shFF49297D;
    weight_mem[1011] = 32'shFF0F5865;
    weight_mem[1012] = 32'sh014D71DC;
    weight_mem[1013] = 32'shFDB3B7B0;
    weight_mem[1014] = 32'shFF5DD5C8;
    weight_mem[1015] = 32'shFF3B8867;
    weight_mem[1016] = 32'shFC0682DC;
    weight_mem[1017] = 32'shFF5B4FA9;
    weight_mem[1018] = 32'shFF6FBD06;
    weight_mem[1019] = 32'shFC4D8184;
    weight_mem[1020] = 32'shFC00C49C;
    weight_mem[1021] = 32'shFFBC04FA;
    weight_mem[1022] = 32'sh02340CAC;
    weight_mem[1023] = 32'sh00B5261B;
    weight_mem[1024] = 32'shFD9F1DFC;
    weight_mem[1025] = 32'sh0298B9BC;
    weight_mem[1026] = 32'shFEE4E294;
    weight_mem[1027] = 32'sh030EB2A0;
    weight_mem[1028] = 32'sh02711A38;
    weight_mem[1029] = 32'shFEFA264C;
    weight_mem[1030] = 32'sh00C499A8;
    weight_mem[1031] = 32'shF9D3BF18;
    weight_mem[1032] = 32'sh02C59874;
    weight_mem[1033] = 32'sh0035E542;
    weight_mem[1034] = 32'shFF0C3C8F;
    weight_mem[1035] = 32'shFE82EEAE;
    weight_mem[1036] = 32'sh029415B0;
    weight_mem[1037] = 32'shFF68AE09;
    weight_mem[1038] = 32'sh03AA2BBC;
    weight_mem[1039] = 32'shFDAE60B8;
    weight_mem[1040] = 32'shFEA22724;
    weight_mem[1041] = 32'sh03BF2620;
    weight_mem[1042] = 32'shFE3CEB92;
    weight_mem[1043] = 32'sh0051B66E;
    weight_mem[1044] = 32'sh01A81C16;
    weight_mem[1045] = 32'shFFE0324E;
    weight_mem[1046] = 32'shFE748D8A;
    weight_mem[1047] = 32'shFFE25E32;
    weight_mem[1048] = 32'shFF07ABE5;
    weight_mem[1049] = 32'shFB3FCBF8;
    weight_mem[1050] = 32'shFFD58BED;
    weight_mem[1051] = 32'shFCF3EC60;
    weight_mem[1052] = 32'shFB896110;
    weight_mem[1053] = 32'shFEFDD9D4;
    weight_mem[1054] = 32'sh0008352A;
    weight_mem[1055] = 32'sh00F93D86;
    weight_mem[1056] = 32'sh005F07EB;
    weight_mem[1057] = 32'shF8F50A10;
    weight_mem[1058] = 32'sh05E9E8B8;
    weight_mem[1059] = 32'sh07A6B9B8;
    weight_mem[1060] = 32'sh047C4DF0;
    weight_mem[1061] = 32'sh0210BA20;
    weight_mem[1062] = 32'shFEF2F7B6;
    weight_mem[1063] = 32'shF9A2C400;
    weight_mem[1064] = 32'sh09318580;
    weight_mem[1065] = 32'sh00281B13;
    weight_mem[1066] = 32'sh03DFD06C;
    weight_mem[1067] = 32'sh032A7F2C;
    weight_mem[1068] = 32'sh02A98F4C;
    weight_mem[1069] = 32'shFA9AD4F0;
    weight_mem[1070] = 32'sh001DBFDE;
    weight_mem[1071] = 32'sh006C37F6;
    weight_mem[1072] = 32'shFDB83FCC;
    weight_mem[1073] = 32'shFFE70DF1;
    weight_mem[1074] = 32'shF77A4360;
    weight_mem[1075] = 32'shFC071154;
    weight_mem[1076] = 32'sh05B41AD0;
    weight_mem[1077] = 32'shF3C7EB20;
    weight_mem[1078] = 32'shFB32D090;
    weight_mem[1079] = 32'sh04545520;
    weight_mem[1080] = 32'shF4D5D720;
    weight_mem[1081] = 32'sh08B41880;
    weight_mem[1082] = 32'shF9C6C030;
    weight_mem[1083] = 32'shF807DD70;
    weight_mem[1084] = 32'shF3485300;
    weight_mem[1085] = 32'sh0671C110;
    weight_mem[1086] = 32'shFF6AB812;
    weight_mem[1087] = 32'sh0140A33C;
    weight_mem[1088] = 32'sh054CD9B8;
    weight_mem[1089] = 32'shFFC93DC1;
    weight_mem[1090] = 32'shFD82456C;
    weight_mem[1091] = 32'shF9D25580;
    weight_mem[1092] = 32'sh024FC2DC;
    weight_mem[1093] = 32'sh03C32258;
    weight_mem[1094] = 32'shFE5D3CCC;
    weight_mem[1095] = 32'sh060DD110;
    weight_mem[1096] = 32'shFF498ED4;
    weight_mem[1097] = 32'shF9D50CB8;
    weight_mem[1098] = 32'sh04244088;
    weight_mem[1099] = 32'shFC8793F8;
    weight_mem[1100] = 32'shFF37CC9D;
    weight_mem[1101] = 32'sh00313F2E;
    weight_mem[1102] = 32'sh06474370;
    weight_mem[1103] = 32'shFEF66536;
    weight_mem[1104] = 32'sh017E83D0;
    weight_mem[1105] = 32'shFB4C7060;
    weight_mem[1106] = 32'shFB23F400;
    weight_mem[1107] = 32'sh02954794;
    weight_mem[1108] = 32'sh054A6FC8;
    weight_mem[1109] = 32'shFFB49F64;
    weight_mem[1110] = 32'shFEE7DB60;
    weight_mem[1111] = 32'sh0341F51C;
    weight_mem[1112] = 32'shFC1C6C40;
    weight_mem[1113] = 32'shFC3CD138;
    weight_mem[1114] = 32'sh03E69428;
    weight_mem[1115] = 32'sh017153D8;
    weight_mem[1116] = 32'shFE138F24;
    weight_mem[1117] = 32'shFF004628;
    weight_mem[1118] = 32'shF931EE08;
    weight_mem[1119] = 32'sh00FB5C13;
    weight_mem[1120] = 32'sh00F1FD32;
    weight_mem[1121] = 32'shFF6ED7A9;
    weight_mem[1122] = 32'shFE4F79D4;
    weight_mem[1123] = 32'shFCAC3E94;
    weight_mem[1124] = 32'shFE423366;
    weight_mem[1125] = 32'sh022BB71C;
    weight_mem[1126] = 32'sh00C54BED;
    weight_mem[1127] = 32'sh06058D10;
    weight_mem[1128] = 32'shFCB03724;
    weight_mem[1129] = 32'shFD730DE8;
    weight_mem[1130] = 32'shFD930B08;
    weight_mem[1131] = 32'shFB442548;
    weight_mem[1132] = 32'sh015FF442;
    weight_mem[1133] = 32'shFF6640AB;
    weight_mem[1134] = 32'shFC9B6DE0;
    weight_mem[1135] = 32'shFF1C6348;
    weight_mem[1136] = 32'sh00D61ACB;
    weight_mem[1137] = 32'shFB2BEDB8;
    weight_mem[1138] = 32'sh017743FA;
    weight_mem[1139] = 32'shFF176D3E;
    weight_mem[1140] = 32'sh036F9F04;
    weight_mem[1141] = 32'shFFC6CD4C;
    weight_mem[1142] = 32'sh00F6C1D0;
    weight_mem[1143] = 32'shFD7EFC7C;
    weight_mem[1144] = 32'sh06B5E030;
    weight_mem[1145] = 32'shFF487DCC;
    weight_mem[1146] = 32'shFE9DCE66;
    weight_mem[1147] = 32'sh02C5AB5C;
    weight_mem[1148] = 32'sh006A5656;
    weight_mem[1149] = 32'shFD8726D4;
    weight_mem[1150] = 32'sh06425A80;
    weight_mem[1151] = 32'sh007A3BCA;
    weight_mem[1152] = 32'shFCEB6AF8;
    weight_mem[1153] = 32'shFCAC8BB0;
    weight_mem[1154] = 32'sh004AE280;
    weight_mem[1155] = 32'shFF2C4F4D;
    weight_mem[1156] = 32'sh001518B0;
    weight_mem[1157] = 32'sh00A13F9B;
    weight_mem[1158] = 32'shFE0372B0;
    weight_mem[1159] = 32'shFE8119E8;
    weight_mem[1160] = 32'shFF49CAF7;
    weight_mem[1161] = 32'shFF13264F;
    weight_mem[1162] = 32'sh0271E348;
    weight_mem[1163] = 32'shFEC40672;
    weight_mem[1164] = 32'shFD2115C0;
    weight_mem[1165] = 32'sh0A20BD90;
    weight_mem[1166] = 32'shFD2E6768;
    weight_mem[1167] = 32'sh05125EF0;
    weight_mem[1168] = 32'shFAAD7490;
    weight_mem[1169] = 32'shFBC3FA88;
    weight_mem[1170] = 32'sh0110D4D6;
    weight_mem[1171] = 32'shFE9FCC4A;
    weight_mem[1172] = 32'sh052286A8;
    weight_mem[1173] = 32'shF73ACE50;
    weight_mem[1174] = 32'shFD58FFFC;
    weight_mem[1175] = 32'sh01B8D092;
    weight_mem[1176] = 32'shFE8F778E;
    weight_mem[1177] = 32'sh010B0720;
    weight_mem[1178] = 32'shF9711958;
    weight_mem[1179] = 32'shFEBEFB00;
    weight_mem[1180] = 32'sh01764BDC;
    weight_mem[1181] = 32'shFF360EC5;
    weight_mem[1182] = 32'sh026CA054;
    weight_mem[1183] = 32'sh0262C940;
    weight_mem[1184] = 32'sh036FE984;
    weight_mem[1185] = 32'sh0457CD50;
    weight_mem[1186] = 32'sh032569C0;
    weight_mem[1187] = 32'shFB153FF0;
    weight_mem[1188] = 32'shFE674FDE;
    weight_mem[1189] = 32'sh035F9F70;
    weight_mem[1190] = 32'sh03C61694;
    weight_mem[1191] = 32'shFBD7BBC0;
    weight_mem[1192] = 32'sh06320C98;
    weight_mem[1193] = 32'shF6E9A2B0;
    weight_mem[1194] = 32'shF80A50F8;
    weight_mem[1195] = 32'sh077618C0;
    weight_mem[1196] = 32'sh0180BD26;
    weight_mem[1197] = 32'sh06E20450;
    weight_mem[1198] = 32'sh08100F10;
    weight_mem[1199] = 32'shF96F5198;
    weight_mem[1200] = 32'sh059516F8;
    weight_mem[1201] = 32'shF839D788;
    weight_mem[1202] = 32'shFA9863A0;
    weight_mem[1203] = 32'shFAD73878;
    weight_mem[1204] = 32'shFAFEC220;
    weight_mem[1205] = 32'shF8CF67A8;
    weight_mem[1206] = 32'sh0491F328;
    weight_mem[1207] = 32'shF89A72C8;
    weight_mem[1208] = 32'sh05605358;
    weight_mem[1209] = 32'sh05E248B8;
    weight_mem[1210] = 32'sh025570E8;
    weight_mem[1211] = 32'sh05EAA1E0;
    weight_mem[1212] = 32'shFF48CD3E;
    weight_mem[1213] = 32'shFE0754B4;
    weight_mem[1214] = 32'shFC0AF134;
    weight_mem[1215] = 32'shFB5A0BD0;
    weight_mem[1216] = 32'shFE9B8F4A;
    weight_mem[1217] = 32'shFC6CCEF4;
    weight_mem[1218] = 32'shFD263548;
    weight_mem[1219] = 32'sh03C6B8CC;
    weight_mem[1220] = 32'sh03F05AD0;
    weight_mem[1221] = 32'sh0124908C;
    weight_mem[1222] = 32'shFD4FF0E4;
    weight_mem[1223] = 32'sh025AC204;
    weight_mem[1224] = 32'shFB23B8B0;
    weight_mem[1225] = 32'sh07866FB8;
    weight_mem[1226] = 32'sh0713CB00;
    weight_mem[1227] = 32'shFB0415C0;
    weight_mem[1228] = 32'shFC1586C4;
    weight_mem[1229] = 32'shF9E25CF8;
    weight_mem[1230] = 32'shF94F83A8;
    weight_mem[1231] = 32'sh057D0AA8;
    weight_mem[1232] = 32'shFBD7ADD0;
    weight_mem[1233] = 32'sh04887048;
    weight_mem[1234] = 32'sh040A3A88;
    weight_mem[1235] = 32'sh04208E70;
    weight_mem[1236] = 32'sh03E82A2C;
    weight_mem[1237] = 32'sh05319298;
    weight_mem[1238] = 32'shFC8050E4;
    weight_mem[1239] = 32'sh068FE470;
    weight_mem[1240] = 32'shFC1C4BD0;
    weight_mem[1241] = 32'shFB4CEB48;
    weight_mem[1242] = 32'shFE355DBE;
    weight_mem[1243] = 32'sh02ED2B5C;
    weight_mem[1244] = 32'shFB5D61A0;
    weight_mem[1245] = 32'sh017CC066;
    weight_mem[1246] = 32'sh030F4AC0;
    weight_mem[1247] = 32'sh04628088;
    weight_mem[1248] = 32'shFB600508;
    weight_mem[1249] = 32'shFBA49490;
    weight_mem[1250] = 32'shFCB4A90C;
    weight_mem[1251] = 32'sh04EA4CC8;
    weight_mem[1252] = 32'sh040EB0D0;
    weight_mem[1253] = 32'shF993D828;
    weight_mem[1254] = 32'shFC47C700;
    weight_mem[1255] = 32'shFCFDF030;
    weight_mem[1256] = 32'shF9B6E4C8;
    weight_mem[1257] = 32'sh09107CA0;
    weight_mem[1258] = 32'sh080DA570;
    weight_mem[1259] = 32'shF8D98C10;
    weight_mem[1260] = 32'shFD3A477C;
    weight_mem[1261] = 32'shF9233EA8;
    weight_mem[1262] = 32'shF7F52420;
    weight_mem[1263] = 32'sh069590E0;
    weight_mem[1264] = 32'shFA796FE0;
    weight_mem[1265] = 32'sh07C2ACA0;
    weight_mem[1266] = 32'sh055A8ED8;
    weight_mem[1267] = 32'sh0529B838;
    weight_mem[1268] = 32'sh050A7CB0;
    weight_mem[1269] = 32'sh07441BB8;
    weight_mem[1270] = 32'shFB5B18B0;
    weight_mem[1271] = 32'sh077E11F8;
    weight_mem[1272] = 32'shFA80C170;
    weight_mem[1273] = 32'shFA03BCF8;
    weight_mem[1274] = 32'shFDB2EE54;
    weight_mem[1275] = 32'sh0185ADAC;
    weight_mem[1276] = 32'shFC886430;
    weight_mem[1277] = 32'sh01F944BE;
    weight_mem[1278] = 32'sh03E774C0;
    weight_mem[1279] = 32'sh03BA78D4;
    weight_mem[1280] = 32'shFF9F7BA0;
    weight_mem[1281] = 32'shFBBF39D8;
    weight_mem[1282] = 32'sh0086A84B;
end

// Pattern B weights
initial begin
    weight_b_mem[   0] = 32'shFFFD87AA;
    weight_b_mem[   1] = 32'sh11102B40;
    weight_b_mem[   2] = 32'sh0B10F560;
    weight_b_mem[   3] = 32'sh00073E6D;
    weight_b_mem[   4] = 32'shE4C52BA0;
    weight_b_mem[   5] = 32'shD0AE5A00;
    weight_b_mem[   6] = 32'shFFF91E4C;
    weight_b_mem[   7] = 32'sh13D084C0;
    weight_b_mem[   8] = 32'sh12E63BC0;
    weight_b_mem[   9] = 32'sh000687E9;
    weight_b_mem[  10] = 32'sh215B9A80;
    weight_b_mem[  11] = 32'shEA0FCC60;
    weight_b_mem[  12] = 32'shFFF6631C;
    weight_b_mem[  13] = 32'sh143CF040;
    weight_b_mem[  14] = 32'sh2EEEE880;
    weight_b_mem[  15] = 32'sh00095BAD;
    weight_b_mem[  16] = 32'sh226F15C0;
    weight_b_mem[  17] = 32'shEC340580;
    weight_b_mem[  18] = 32'sh00018EE7;
    weight_b_mem[  19] = 32'shE72D7500;
    weight_b_mem[  20] = 32'shFBE07C98;
    weight_b_mem[  21] = 32'sh0008D586;
    weight_b_mem[  22] = 32'sh0A67C970;
    weight_b_mem[  23] = 32'shD6725700;
    weight_b_mem[  24] = 32'shFFF66201;
    weight_b_mem[  25] = 32'sh00E045FE;
    weight_b_mem[  26] = 32'sh27AC0200;
    weight_b_mem[  27] = 32'shFFFCF9CE;
    weight_b_mem[  28] = 32'shFF428320;
    weight_b_mem[  29] = 32'sh0B45C540;
    weight_b_mem[  30] = 32'shFFF4A482;
    weight_b_mem[  31] = 32'shF260F030;
    weight_b_mem[  32] = 32'sh2B110540;
    weight_b_mem[  33] = 32'shFFFFA69B;
    weight_b_mem[  34] = 32'shF129B820;
    weight_b_mem[  35] = 32'shFB900410;
    weight_b_mem[  36] = 32'shFFFDE156;
    weight_b_mem[  37] = 32'shF8D014C8;
    weight_b_mem[  38] = 32'sh18F2DEC0;
    weight_b_mem[  39] = 32'sh000BE102;
    weight_b_mem[  40] = 32'sh20C661C0;
    weight_b_mem[  41] = 32'sh164A3760;
    weight_b_mem[  42] = 32'sh0000FCF8;
    weight_b_mem[  43] = 32'shED064800;
    weight_b_mem[  44] = 32'shF60C6470;
    weight_b_mem[  45] = 32'shFFFBF5E2;
    weight_b_mem[  46] = 32'shF7FDBD30;
    weight_b_mem[  47] = 32'sh0F47D050;
    weight_b_mem[  48] = 32'sh00013BAC;
    weight_b_mem[  49] = 32'shF9CBBA90;
    weight_b_mem[  50] = 32'shE6D9CB80;
    weight_b_mem[  51] = 32'sh00067FA8;
    weight_b_mem[  52] = 32'sh178895E0;
    weight_b_mem[  53] = 32'shEDCEDE00;
    weight_b_mem[  54] = 32'shFFFC7CBA;
    weight_b_mem[  55] = 32'shE69DBCE0;
    weight_b_mem[  56] = 32'sh15B00AA0;
    weight_b_mem[  57] = 32'shFFF76293;
    weight_b_mem[  58] = 32'shEEA83180;
    weight_b_mem[  59] = 32'sh2B89DAC0;
    weight_b_mem[  60] = 32'shFFFCB9F9;
    weight_b_mem[  61] = 32'shF3D9B740;
    weight_b_mem[  62] = 32'sh09694AE0;
    weight_b_mem[  63] = 32'sh0004DCD7;
    weight_b_mem[  64] = 32'sh10D03D60;
    weight_b_mem[  65] = 32'shF8F61820;
    weight_b_mem[  66] = 32'shFFFE03FA;
    weight_b_mem[  67] = 32'sh0CAC4790;
    weight_b_mem[  68] = 32'shFE97E8CE;
    weight_b_mem[  69] = 32'sh0004E40B;
    weight_b_mem[  70] = 32'shFD7D6000;
    weight_b_mem[  71] = 32'shDE8249C0;
    weight_b_mem[  72] = 32'sh00012F03;
    weight_b_mem[  73] = 32'shD64F4640;
    weight_b_mem[  74] = 32'shF78D5D40;
    weight_b_mem[  75] = 32'shFFFE76E2;
    weight_b_mem[  76] = 32'sh2C666F00;
    weight_b_mem[  77] = 32'sh0125B19E;
    weight_b_mem[  78] = 32'shFFF74A80;
    weight_b_mem[  79] = 32'sh03F95D10;
    weight_b_mem[  80] = 32'sh1CEA8240;
    weight_b_mem[  81] = 32'shFFFDB5E4;
    weight_b_mem[  82] = 32'shD5B84480;
    weight_b_mem[  83] = 32'sh05F65AB8;
    weight_b_mem[  84] = 32'shFFFF209E;
    weight_b_mem[  85] = 32'shD6E09A40;
    weight_b_mem[  86] = 32'shEABEDF20;
    weight_b_mem[  87] = 32'shFFF6387E;
    weight_b_mem[  88] = 32'shEB2D3AC0;
    weight_b_mem[  89] = 32'sh27401B00;
    weight_b_mem[  90] = 32'shFFFD2084;
    weight_b_mem[  91] = 32'sh069DC4C0;
    weight_b_mem[  92] = 32'sh05AA3168;
    weight_b_mem[  93] = 32'sh0009D23E;
    weight_b_mem[  94] = 32'sh0E5716E0;
    weight_b_mem[  95] = 32'shDA273D00;
    weight_b_mem[  96] = 32'sh51B95E00;
    weight_b_mem[  97] = 32'shC4007980;
    weight_b_mem[  98] = 32'sh26E0FD80;
    weight_b_mem[  99] = 32'shB0750100;
    weight_b_mem[ 100] = 32'sh40BC3F80;
    weight_b_mem[ 101] = 32'sh3A97DCC0;
    weight_b_mem[ 102] = 32'sh2A91C880;
    weight_b_mem[ 103] = 32'sh0447A048;
    weight_b_mem[ 104] = 32'sh00F608B1;
    weight_b_mem[ 105] = 32'sh351ADA40;
    weight_b_mem[ 106] = 32'sh5AB93980;
    weight_b_mem[ 107] = 32'shE1F7EA40;
    weight_b_mem[ 108] = 32'shF3E16980;
    weight_b_mem[ 109] = 32'shF4589380;
    weight_b_mem[ 110] = 32'sh20491800;
    weight_b_mem[ 111] = 32'sh3B3E7580;
    weight_b_mem[ 112] = 32'sh4288CE00;
    weight_b_mem[ 113] = 32'sh086B6810;
    weight_b_mem[ 114] = 32'shD0196E00;
    weight_b_mem[ 115] = 32'shBE306C80;
    weight_b_mem[ 116] = 32'shEDB424C0;
    weight_b_mem[ 117] = 32'sh4DAAA880;
    weight_b_mem[ 118] = 32'sh0F74BBE0;
    weight_b_mem[ 119] = 32'sh07F99EF0;
    weight_b_mem[ 120] = 32'sh38634640;
    weight_b_mem[ 121] = 32'shF6DD52A0;
    weight_b_mem[ 122] = 32'sh653BE080;
    weight_b_mem[ 123] = 32'sh3D4B2580;
    weight_b_mem[ 124] = 32'shD4027C40;
    weight_b_mem[ 125] = 32'sh0DAA34C0;
    weight_b_mem[ 126] = 32'sh5B281300;
    weight_b_mem[ 127] = 32'sh516EC100;
    weight_b_mem[ 128] = 32'sh07E527A0;
    weight_b_mem[ 129] = 32'shFD691FC0;
    weight_b_mem[ 130] = 32'shF54924B0;
    weight_b_mem[ 131] = 32'sh007DF581;
    weight_b_mem[ 132] = 32'shFC7CD82C;
    weight_b_mem[ 133] = 32'shFB9F8FC8;
    weight_b_mem[ 134] = 32'sh00E0F4E5;
    weight_b_mem[ 135] = 32'shFF64B74A;
    weight_b_mem[ 136] = 32'shFE70778E;
    weight_b_mem[ 137] = 32'shFCCC3358;
    weight_b_mem[ 138] = 32'shFEF6BD92;
    weight_b_mem[ 139] = 32'sh04E67620;
    weight_b_mem[ 140] = 32'sh01B68648;
    weight_b_mem[ 141] = 32'sh01769BF4;
    weight_b_mem[ 142] = 32'sh0083831D;
    weight_b_mem[ 143] = 32'shFC12ECC4;
    weight_b_mem[ 144] = 32'shFC9E3668;
    weight_b_mem[ 145] = 32'shFC9DB57C;
    weight_b_mem[ 146] = 32'shFE2D73D8;
    weight_b_mem[ 147] = 32'shFBC86230;
    weight_b_mem[ 148] = 32'shFC5332B4;
    weight_b_mem[ 149] = 32'sh04875F70;
    weight_b_mem[ 150] = 32'shFB742058;
    weight_b_mem[ 151] = 32'sh02164D14;
    weight_b_mem[ 152] = 32'shF81374E8;
    weight_b_mem[ 153] = 32'sh06B018E0;
    weight_b_mem[ 154] = 32'sh0067C29B;
    weight_b_mem[ 155] = 32'shF60E33E0;
    weight_b_mem[ 156] = 32'sh00887964;
    weight_b_mem[ 157] = 32'shFBFE3F48;
    weight_b_mem[ 158] = 32'shFD6A7EEC;
    weight_b_mem[ 159] = 32'shFFC01DF1;
    weight_b_mem[ 160] = 32'shFD42276C;
    weight_b_mem[ 161] = 32'sh013195F4;
    weight_b_mem[ 162] = 32'sh03CEE814;
    weight_b_mem[ 163] = 32'shFE0BDC0E;
    weight_b_mem[ 164] = 32'sh00938738;
    weight_b_mem[ 165] = 32'shFDB3ADF4;
    weight_b_mem[ 166] = 32'sh085BF8C0;
    weight_b_mem[ 167] = 32'sh02574E14;
    weight_b_mem[ 168] = 32'shFF8242CA;
    weight_b_mem[ 169] = 32'shFEE5619C;
    weight_b_mem[ 170] = 32'sh01101AFE;
    weight_b_mem[ 171] = 32'shFBB3B100;
    weight_b_mem[ 172] = 32'sh065E8588;
    weight_b_mem[ 173] = 32'shFFB3E2C0;
    weight_b_mem[ 174] = 32'shFAD298F0;
    weight_b_mem[ 175] = 32'shFFE1B727;
    weight_b_mem[ 176] = 32'sh020B9128;
    weight_b_mem[ 177] = 32'sh05E8EB10;
    weight_b_mem[ 178] = 32'shFE1073A4;
    weight_b_mem[ 179] = 32'sh0082ADEB;
    weight_b_mem[ 180] = 32'sh007C6C7A;
    weight_b_mem[ 181] = 32'shFA54C030;
    weight_b_mem[ 182] = 32'shFB9E96F0;
    weight_b_mem[ 183] = 32'shFBE2B7A0;
    weight_b_mem[ 184] = 32'sh02B368A8;
    weight_b_mem[ 185] = 32'shFDC2D940;
    weight_b_mem[ 186] = 32'sh00309702;
    weight_b_mem[ 187] = 32'shFD3E5B40;
    weight_b_mem[ 188] = 32'sh039D8D8C;
    weight_b_mem[ 189] = 32'sh007040D0;
    weight_b_mem[ 190] = 32'sh0468B308;
    weight_b_mem[ 191] = 32'shFDB52458;
    weight_b_mem[ 192] = 32'shF6E30D00;
    weight_b_mem[ 193] = 32'shF9CF4E98;
    weight_b_mem[ 194] = 32'shFDE8ACFC;
    weight_b_mem[ 195] = 32'shFACDC7C0;
    weight_b_mem[ 196] = 32'shFB4D8138;
    weight_b_mem[ 197] = 32'shFC753F10;
    weight_b_mem[ 198] = 32'sh081B89C0;
    weight_b_mem[ 199] = 32'sh027D5058;
    weight_b_mem[ 200] = 32'sh004344DA;
    weight_b_mem[ 201] = 32'sh028913D4;
    weight_b_mem[ 202] = 32'sh017ED1EA;
    weight_b_mem[ 203] = 32'sh0508ACE8;
    weight_b_mem[ 204] = 32'sh000995AC;
    weight_b_mem[ 205] = 32'shFE71ACD4;
    weight_b_mem[ 206] = 32'sh06195678;
    weight_b_mem[ 207] = 32'shFCFCAA8C;
    weight_b_mem[ 208] = 32'sh010AE9F8;
    weight_b_mem[ 209] = 32'sh028219F8;
    weight_b_mem[ 210] = 32'sh03ACFFDC;
    weight_b_mem[ 211] = 32'shFBA54EC8;
    weight_b_mem[ 212] = 32'sh0071E9EA;
    weight_b_mem[ 213] = 32'shFD613594;
    weight_b_mem[ 214] = 32'sh07EB91B8;
    weight_b_mem[ 215] = 32'sh02812790;
    weight_b_mem[ 216] = 32'sh05D342B0;
    weight_b_mem[ 217] = 32'shF9D060C0;
    weight_b_mem[ 218] = 32'sh03B462E0;
    weight_b_mem[ 219] = 32'sh0F2CACD0;
    weight_b_mem[ 220] = 32'sh02A1C244;
    weight_b_mem[ 221] = 32'sh02961208;
    weight_b_mem[ 222] = 32'sh06723CB0;
    weight_b_mem[ 223] = 32'sh02ADB120;
    weight_b_mem[ 224] = 32'sh0188ADF4;
    weight_b_mem[ 225] = 32'shFC1C9E84;
    weight_b_mem[ 226] = 32'sh05553B78;
    weight_b_mem[ 227] = 32'sh07936FB0;
    weight_b_mem[ 228] = 32'shFB9B9D78;
    weight_b_mem[ 229] = 32'sh0471BF40;
    weight_b_mem[ 230] = 32'shFB46BA80;
    weight_b_mem[ 231] = 32'sh02A99600;
    weight_b_mem[ 232] = 32'shFC642C3C;
    weight_b_mem[ 233] = 32'shFC24A228;
    weight_b_mem[ 234] = 32'shFF5DAA66;
    weight_b_mem[ 235] = 32'shFD5D4458;
    weight_b_mem[ 236] = 32'shFCE895FC;
    weight_b_mem[ 237] = 32'sh021083EC;
    weight_b_mem[ 238] = 32'shFEB61F22;
    weight_b_mem[ 239] = 32'shF9DDD098;
    weight_b_mem[ 240] = 32'shFFB930B2;
    weight_b_mem[ 241] = 32'shFC0146C0;
    weight_b_mem[ 242] = 32'shFCF41310;
    weight_b_mem[ 243] = 32'sh048463C0;
    weight_b_mem[ 244] = 32'shFFE22D89;
    weight_b_mem[ 245] = 32'sh054CA808;
    weight_b_mem[ 246] = 32'sh05795F48;
    weight_b_mem[ 247] = 32'sh069CBF78;
    weight_b_mem[ 248] = 32'sh015B77E2;
    weight_b_mem[ 249] = 32'shFB77E9D8;
    weight_b_mem[ 250] = 32'shFDFD31F4;
    weight_b_mem[ 251] = 32'sh04052778;
    weight_b_mem[ 252] = 32'sh0094D5DD;
    weight_b_mem[ 253] = 32'sh04786E78;
    weight_b_mem[ 254] = 32'shFE9FBB96;
    weight_b_mem[ 255] = 32'shFF58FA76;
    weight_b_mem[ 256] = 32'sh03189A20;
    weight_b_mem[ 257] = 32'sh00823D11;
    weight_b_mem[ 258] = 32'sh01FFE462;
    weight_b_mem[ 259] = 32'sh01B3D8C6;
    weight_b_mem[ 260] = 32'sh0213310C;
    weight_b_mem[ 261] = 32'sh05461258;
    weight_b_mem[ 262] = 32'sh0191AF20;
    weight_b_mem[ 263] = 32'sh023993E0;
    weight_b_mem[ 264] = 32'sh006043A2;
    weight_b_mem[ 265] = 32'shF98430C8;
    weight_b_mem[ 266] = 32'shFE4F7E1E;
    weight_b_mem[ 267] = 32'shFAF24460;
    weight_b_mem[ 268] = 32'sh00A1597F;
    weight_b_mem[ 269] = 32'sh0493A0C8;
    weight_b_mem[ 270] = 32'shFC4F2898;
    weight_b_mem[ 271] = 32'shFC346F18;
    weight_b_mem[ 272] = 32'sh01471968;
    weight_b_mem[ 273] = 32'sh0031534E;
    weight_b_mem[ 274] = 32'sh045B4D60;
    weight_b_mem[ 275] = 32'shFDC63408;
    weight_b_mem[ 276] = 32'sh03F67328;
    weight_b_mem[ 277] = 32'sh02E24B88;
    weight_b_mem[ 278] = 32'shFC005924;
    weight_b_mem[ 279] = 32'shFC57D3F4;
    weight_b_mem[ 280] = 32'sh0474CB38;
    weight_b_mem[ 281] = 32'sh01D74BB8;
    weight_b_mem[ 282] = 32'sh06292CF0;
    weight_b_mem[ 283] = 32'sh03DF1704;
    weight_b_mem[ 284] = 32'shFEDB6052;
    weight_b_mem[ 285] = 32'sh042DAB20;
    weight_b_mem[ 286] = 32'shFC524B38;
    weight_b_mem[ 287] = 32'sh01F937CA;
    weight_b_mem[ 288] = 32'shFB2BC130;
    weight_b_mem[ 289] = 32'sh00C84F5E;
    weight_b_mem[ 290] = 32'shFC829A10;
    weight_b_mem[ 291] = 32'shFC9C8D7C;
    weight_b_mem[ 292] = 32'shFF55E4A3;
    weight_b_mem[ 293] = 32'sh0040AC26;
    weight_b_mem[ 294] = 32'shFB6AF4B0;
    weight_b_mem[ 295] = 32'shFA38E880;
    weight_b_mem[ 296] = 32'sh0A706020;
    weight_b_mem[ 297] = 32'sh070BF600;
    weight_b_mem[ 298] = 32'shFD59B940;
    weight_b_mem[ 299] = 32'shFC586A84;
    weight_b_mem[ 300] = 32'sh02B79684;
    weight_b_mem[ 301] = 32'sh05D2D908;
    weight_b_mem[ 302] = 32'sh02336518;
    weight_b_mem[ 303] = 32'sh0667EA68;
    weight_b_mem[ 304] = 32'shFE202F5A;
    weight_b_mem[ 305] = 32'sh034EAA90;
    weight_b_mem[ 306] = 32'shFED46D2E;
    weight_b_mem[ 307] = 32'shFFE5DFAB;
    weight_b_mem[ 308] = 32'shFDF52F7C;
    weight_b_mem[ 309] = 32'shFFCA99F3;
    weight_b_mem[ 310] = 32'shFF044DC7;
    weight_b_mem[ 311] = 32'shFB72F348;
    weight_b_mem[ 312] = 32'sh03E3980C;
    weight_b_mem[ 313] = 32'sh020EAF1C;
    weight_b_mem[ 314] = 32'sh07D0DC00;
    weight_b_mem[ 315] = 32'shFAB7A270;
    weight_b_mem[ 316] = 32'shFBE5F098;
    weight_b_mem[ 317] = 32'shFDF40890;
    weight_b_mem[ 318] = 32'shFF3703A5;
    weight_b_mem[ 319] = 32'shFEC2963C;
    weight_b_mem[ 320] = 32'sh01C280E2;
    weight_b_mem[ 321] = 32'shFAD047B0;
    weight_b_mem[ 322] = 32'sh02C9D040;
    weight_b_mem[ 323] = 32'shFE2CBD02;
    weight_b_mem[ 324] = 32'shFB0E19F0;
    weight_b_mem[ 325] = 32'shFF3F927C;
    weight_b_mem[ 326] = 32'sh0B3178C0;
    weight_b_mem[ 327] = 32'shF9D9C838;
    weight_b_mem[ 328] = 32'sh06194C10;
    weight_b_mem[ 329] = 32'sh003B6F0A;
    weight_b_mem[ 330] = 32'sh002D890B;
    weight_b_mem[ 331] = 32'sh02AB2270;
    weight_b_mem[ 332] = 32'shFB179DB8;
    weight_b_mem[ 333] = 32'shFDC407E0;
    weight_b_mem[ 334] = 32'sh014FCBCE;
    weight_b_mem[ 335] = 32'shFEF0E06C;
    weight_b_mem[ 336] = 32'sh02E4B934;
    weight_b_mem[ 337] = 32'sh05295178;
    weight_b_mem[ 338] = 32'shFDB3FA58;
    weight_b_mem[ 339] = 32'sh02FC0B2C;
    weight_b_mem[ 340] = 32'shFEB30062;
    weight_b_mem[ 341] = 32'sh00163465;
    weight_b_mem[ 342] = 32'sh04CD9FC8;
    weight_b_mem[ 343] = 32'shFC909ED8;
    weight_b_mem[ 344] = 32'shF8B47E00;
    weight_b_mem[ 345] = 32'shF828FF60;
    weight_b_mem[ 346] = 32'sh04ECAC78;
    weight_b_mem[ 347] = 32'sh07208C48;
    weight_b_mem[ 348] = 32'shFF84781A;
    weight_b_mem[ 349] = 32'sh00E7FC38;
    weight_b_mem[ 350] = 32'shF8559B58;
    weight_b_mem[ 351] = 32'sh0426E950;
    weight_b_mem[ 352] = 32'sh06E10B60;
    weight_b_mem[ 353] = 32'shFF941277;
    weight_b_mem[ 354] = 32'sh0320CFA8;
    weight_b_mem[ 355] = 32'shFEA83E5A;
    weight_b_mem[ 356] = 32'shFEE7B442;
    weight_b_mem[ 357] = 32'shFABD4918;
    weight_b_mem[ 358] = 32'shFC187498;
    weight_b_mem[ 359] = 32'shFC0CFFC8;
    weight_b_mem[ 360] = 32'shFE4C03CA;
    weight_b_mem[ 361] = 32'shFC5F9C20;
    weight_b_mem[ 362] = 32'shFDA91DFC;
    weight_b_mem[ 363] = 32'sh02E92A34;
    weight_b_mem[ 364] = 32'sh06ACDE18;
    weight_b_mem[ 365] = 32'sh013E6A80;
    weight_b_mem[ 366] = 32'sh04AF0F50;
    weight_b_mem[ 367] = 32'sh06533F10;
    weight_b_mem[ 368] = 32'shFDD21DD0;
    weight_b_mem[ 369] = 32'shFD9D80C4;
    weight_b_mem[ 370] = 32'shFDF6FA20;
    weight_b_mem[ 371] = 32'sh01998F4E;
    weight_b_mem[ 372] = 32'shFE5ED80E;
    weight_b_mem[ 373] = 32'shFB547D90;
    weight_b_mem[ 374] = 32'shFDE3CEF4;
    weight_b_mem[ 375] = 32'shFA488870;
    weight_b_mem[ 376] = 32'sh06605A48;
    weight_b_mem[ 377] = 32'sh000D9818;
    weight_b_mem[ 378] = 32'shFFB89598;
    weight_b_mem[ 379] = 32'shFE082D8A;
    weight_b_mem[ 380] = 32'sh03CB64C4;
    weight_b_mem[ 381] = 32'sh02C86278;
    weight_b_mem[ 382] = 32'sh04363D20;
    weight_b_mem[ 383] = 32'shFE4A08D4;
    weight_b_mem[ 384] = 32'sh01588574;
    weight_b_mem[ 385] = 32'sh02D6BEE0;
    weight_b_mem[ 386] = 32'shFF0D5719;
    weight_b_mem[ 387] = 32'shFD59B970;
    weight_b_mem[ 388] = 32'sh03D08850;
    weight_b_mem[ 389] = 32'shFCD51D24;
    weight_b_mem[ 390] = 32'sh020FAF48;
    weight_b_mem[ 391] = 32'shFDE12230;
    weight_b_mem[ 392] = 32'shFBEFABF8;
    weight_b_mem[ 393] = 32'shFC25226C;
    weight_b_mem[ 394] = 32'sh00ADA3D6;
    weight_b_mem[ 395] = 32'shFC831900;
    weight_b_mem[ 396] = 32'shFC17E27C;
    weight_b_mem[ 397] = 32'sh03E77DC8;
    weight_b_mem[ 398] = 32'sh001BEBF6;
    weight_b_mem[ 399] = 32'sh011ACF44;
    weight_b_mem[ 400] = 32'sh03EA45D4;
    weight_b_mem[ 401] = 32'shFF3096F0;
    weight_b_mem[ 402] = 32'sh0367C26C;
    weight_b_mem[ 403] = 32'shFF4AADCA;
    weight_b_mem[ 404] = 32'sh075CB688;
    weight_b_mem[ 405] = 32'sh02EB99FC;
    weight_b_mem[ 406] = 32'shFAE38EC0;
    weight_b_mem[ 407] = 32'sh00F36986;
    weight_b_mem[ 408] = 32'shF6B0C7C0;
    weight_b_mem[ 409] = 32'shFD6F7F98;
    weight_b_mem[ 410] = 32'shFF0892E3;
    weight_b_mem[ 411] = 32'sh059D2900;
    weight_b_mem[ 412] = 32'shFEA458B0;
    weight_b_mem[ 413] = 32'shFDCD06FC;
    weight_b_mem[ 414] = 32'shFC4FF394;
    weight_b_mem[ 415] = 32'sh02FE6E60;
    weight_b_mem[ 416] = 32'sh05432608;
    weight_b_mem[ 417] = 32'shFF3703D6;
    weight_b_mem[ 418] = 32'sh03C3B31C;
    weight_b_mem[ 419] = 32'shFDA026D0;
    weight_b_mem[ 420] = 32'sh0053494C;
    weight_b_mem[ 421] = 32'shFC609C8C;
    weight_b_mem[ 422] = 32'sh04C3C540;
    weight_b_mem[ 423] = 32'shFB14A2D8;
    weight_b_mem[ 424] = 32'shF9BCAAE0;
    weight_b_mem[ 425] = 32'shFC78C28C;
    weight_b_mem[ 426] = 32'sh02B44508;
    weight_b_mem[ 427] = 32'sh04CD0C70;
    weight_b_mem[ 428] = 32'sh051177F8;
    weight_b_mem[ 429] = 32'sh01C82A2A;
    weight_b_mem[ 430] = 32'shFD9CCC50;
    weight_b_mem[ 431] = 32'shFDC821F0;
    weight_b_mem[ 432] = 32'shFA161ED8;
    weight_b_mem[ 433] = 32'sh06A95A48;
    weight_b_mem[ 434] = 32'shFC77E2EC;
    weight_b_mem[ 435] = 32'sh026AE848;
    weight_b_mem[ 436] = 32'shF5EBE5D0;
    weight_b_mem[ 437] = 32'sh09AB85F0;
    weight_b_mem[ 438] = 32'sh03A902DC;
    weight_b_mem[ 439] = 32'sh02006590;
    weight_b_mem[ 440] = 32'shF368DA20;
    weight_b_mem[ 441] = 32'sh0261E4D4;
    weight_b_mem[ 442] = 32'shF6B9C690;
    weight_b_mem[ 443] = 32'shFE3D9FB6;
    weight_b_mem[ 444] = 32'sh05043F48;
    weight_b_mem[ 445] = 32'shFFD76505;
    weight_b_mem[ 446] = 32'sh01ED9180;
    weight_b_mem[ 447] = 32'sh031F5BD4;
    weight_b_mem[ 448] = 32'sh05290908;
    weight_b_mem[ 449] = 32'shFC8AC8E8;
    weight_b_mem[ 450] = 32'sh048DBB80;
    weight_b_mem[ 451] = 32'sh00527636;
    weight_b_mem[ 452] = 32'shFD955CC4;
    weight_b_mem[ 453] = 32'sh023982C0;
    weight_b_mem[ 454] = 32'shF97A8640;
    weight_b_mem[ 455] = 32'sh01F7BEFA;
    weight_b_mem[ 456] = 32'shFC3472B4;
    weight_b_mem[ 457] = 32'sh02C894A8;
    weight_b_mem[ 458] = 32'sh02866CC0;
    weight_b_mem[ 459] = 32'shFB5B9B88;
    weight_b_mem[ 460] = 32'shFC6FB9AC;
    weight_b_mem[ 461] = 32'shFAA850C0;
    weight_b_mem[ 462] = 32'shFB727830;
    weight_b_mem[ 463] = 32'shFF202682;
    weight_b_mem[ 464] = 32'sh06ED55E8;
    weight_b_mem[ 465] = 32'shFE1D53EC;
    weight_b_mem[ 466] = 32'sh0091B457;
    weight_b_mem[ 467] = 32'shFEEA57B8;
    weight_b_mem[ 468] = 32'shFFCF150B;
    weight_b_mem[ 469] = 32'sh02781534;
    weight_b_mem[ 470] = 32'sh011A8932;
    weight_b_mem[ 471] = 32'shFBBB2A48;
    weight_b_mem[ 472] = 32'shFC68C4F8;
    weight_b_mem[ 473] = 32'sh0086CB64;
    weight_b_mem[ 474] = 32'shFBF68300;
    weight_b_mem[ 475] = 32'shFD596018;
    weight_b_mem[ 476] = 32'sh00B31FB4;
    weight_b_mem[ 477] = 32'sh02456EEC;
    weight_b_mem[ 478] = 32'sh06BB2D88;
    weight_b_mem[ 479] = 32'sh01BE2AA0;
    weight_b_mem[ 480] = 32'sh00CF777F;
    weight_b_mem[ 481] = 32'sh00D4EB76;
    weight_b_mem[ 482] = 32'shFD3DB750;
    weight_b_mem[ 483] = 32'shFFD93730;
    weight_b_mem[ 484] = 32'sh0090E946;
    weight_b_mem[ 485] = 32'shFC51EDBC;
    weight_b_mem[ 486] = 32'sh068F8840;
    weight_b_mem[ 487] = 32'sh03D9F9B0;
    weight_b_mem[ 488] = 32'sh019D43D2;
    weight_b_mem[ 489] = 32'shFB7E4A78;
    weight_b_mem[ 490] = 32'shFE873222;
    weight_b_mem[ 491] = 32'sh0313650C;
    weight_b_mem[ 492] = 32'sh04AB6738;
    weight_b_mem[ 493] = 32'shFDD4BB84;
    weight_b_mem[ 494] = 32'shFFA74F5C;
    weight_b_mem[ 495] = 32'sh0324B6A8;
    weight_b_mem[ 496] = 32'sh003D4BC4;
    weight_b_mem[ 497] = 32'sh01CE812E;
    weight_b_mem[ 498] = 32'shFC178180;
    weight_b_mem[ 499] = 32'shFB1A2668;
    weight_b_mem[ 500] = 32'sh05D3FF80;
    weight_b_mem[ 501] = 32'sh01F79200;
    weight_b_mem[ 502] = 32'shFBE1BB70;
    weight_b_mem[ 503] = 32'shF8E97E38;
    weight_b_mem[ 504] = 32'shF9712550;
    weight_b_mem[ 505] = 32'sh02AF3890;
    weight_b_mem[ 506] = 32'sh0399DDC8;
    weight_b_mem[ 507] = 32'shF9DFE630;
    weight_b_mem[ 508] = 32'sh03F38DD8;
    weight_b_mem[ 509] = 32'shFBF9B048;
    weight_b_mem[ 510] = 32'shFA7168C8;
    weight_b_mem[ 511] = 32'shFD878ECC;
    weight_b_mem[ 512] = 32'shEF1F3940;
    weight_b_mem[ 513] = 32'sh01EAA7FE;
    weight_b_mem[ 514] = 32'shFBA15080;
    weight_b_mem[ 515] = 32'sh0168E440;
    weight_b_mem[ 516] = 32'sh0312D6F4;
    weight_b_mem[ 517] = 32'sh07989190;
    weight_b_mem[ 518] = 32'shF24E1DF0;
    weight_b_mem[ 519] = 32'shFDFEF230;
    weight_b_mem[ 520] = 32'shFF1F7C84;
    weight_b_mem[ 521] = 32'sh02260728;
    weight_b_mem[ 522] = 32'shF9983270;
    weight_b_mem[ 523] = 32'sh0B7FF350;
    weight_b_mem[ 524] = 32'shFEF53ED4;
    weight_b_mem[ 525] = 32'shFCC30AC0;
    weight_b_mem[ 526] = 32'sh080ED470;
    weight_b_mem[ 527] = 32'sh06F00648;
    weight_b_mem[ 528] = 32'sh012872D6;
    weight_b_mem[ 529] = 32'shF9B6A2D8;
    weight_b_mem[ 530] = 32'sh06C21C30;
    weight_b_mem[ 531] = 32'shFEBBA1F0;
    weight_b_mem[ 532] = 32'sh09BF1110;
    weight_b_mem[ 533] = 32'shF4052EC0;
    weight_b_mem[ 534] = 32'sh0D89B050;
    weight_b_mem[ 535] = 32'sh01A0C1F4;
    weight_b_mem[ 536] = 32'sh0CF4E360;
    weight_b_mem[ 537] = 32'shEC9C4B40;
    weight_b_mem[ 538] = 32'sh032C5E24;
    weight_b_mem[ 539] = 32'sh0FC5AFB0;
    weight_b_mem[ 540] = 32'shFF660887;
    weight_b_mem[ 541] = 32'sh060B6AD0;
    weight_b_mem[ 542] = 32'sh043F22A8;
    weight_b_mem[ 543] = 32'sh007A2A3C;
    weight_b_mem[ 544] = 32'sh0421BA08;
    weight_b_mem[ 545] = 32'sh00442AFE;
    weight_b_mem[ 546] = 32'shF9D05608;
    weight_b_mem[ 547] = 32'shFBCD37D0;
    weight_b_mem[ 548] = 32'sh00730373;
    weight_b_mem[ 549] = 32'shFC9C2848;
    weight_b_mem[ 550] = 32'sh009F98C0;
    weight_b_mem[ 551] = 32'sh067FE190;
    weight_b_mem[ 552] = 32'sh018BD9C0;
    weight_b_mem[ 553] = 32'shF9AE7020;
    weight_b_mem[ 554] = 32'shFC836078;
    weight_b_mem[ 555] = 32'shFAA49F98;
    weight_b_mem[ 556] = 32'shFF1BEF14;
    weight_b_mem[ 557] = 32'shFE5FDB34;
    weight_b_mem[ 558] = 32'shFC3D9840;
    weight_b_mem[ 559] = 32'sh053C08E0;
    weight_b_mem[ 560] = 32'shFE7E617A;
    weight_b_mem[ 561] = 32'sh046D5528;
    weight_b_mem[ 562] = 32'sh0044122A;
    weight_b_mem[ 563] = 32'shFBE8F148;
    weight_b_mem[ 564] = 32'shF8848158;
    weight_b_mem[ 565] = 32'shFFA0AC9A;
    weight_b_mem[ 566] = 32'sh01124E10;
    weight_b_mem[ 567] = 32'shFF645348;
    weight_b_mem[ 568] = 32'sh02D1BD10;
    weight_b_mem[ 569] = 32'shFAC3C3F0;
    weight_b_mem[ 570] = 32'shFDBDA38C;
    weight_b_mem[ 571] = 32'shFEB9BA42;
    weight_b_mem[ 572] = 32'shFC7BAECC;
    weight_b_mem[ 573] = 32'shFE83C7D4;
    weight_b_mem[ 574] = 32'shFA8EEDB0;
    weight_b_mem[ 575] = 32'shFE1E3F64;
    weight_b_mem[ 576] = 32'shFDBBCCEC;
    weight_b_mem[ 577] = 32'sh04B6F3F8;
    weight_b_mem[ 578] = 32'sh056CB9E0;
    weight_b_mem[ 579] = 32'sh03F41940;
    weight_b_mem[ 580] = 32'sh05531378;
    weight_b_mem[ 581] = 32'shFBF1CDF0;
    weight_b_mem[ 582] = 32'sh01B2731E;
    weight_b_mem[ 583] = 32'shFF291CC7;
    weight_b_mem[ 584] = 32'shFC1967C8;
    weight_b_mem[ 585] = 32'shFD50F708;
    weight_b_mem[ 586] = 32'shFA5C11C0;
    weight_b_mem[ 587] = 32'shFB40BCF8;
    weight_b_mem[ 588] = 32'sh024F0234;
    weight_b_mem[ 589] = 32'shFDA422B8;
    weight_b_mem[ 590] = 32'sh056CF730;
    weight_b_mem[ 591] = 32'sh00296433;
    weight_b_mem[ 592] = 32'sh04C7AC08;
    weight_b_mem[ 593] = 32'shFF413224;
    weight_b_mem[ 594] = 32'sh00E46395;
    weight_b_mem[ 595] = 32'shFC3CDCA8;
    weight_b_mem[ 596] = 32'sh008C47AE;
    weight_b_mem[ 597] = 32'shFA7F6AD8;
    weight_b_mem[ 598] = 32'sh072800E0;
    weight_b_mem[ 599] = 32'sh00A1FF0A;
    weight_b_mem[ 600] = 32'sh0A7921F0;
    weight_b_mem[ 601] = 32'shF80B3E60;
    weight_b_mem[ 602] = 32'sh0006417B;
    weight_b_mem[ 603] = 32'sh097C3000;
    weight_b_mem[ 604] = 32'sh084A2B40;
    weight_b_mem[ 605] = 32'shFCE792F8;
    weight_b_mem[ 606] = 32'sh006CE9E6;
    weight_b_mem[ 607] = 32'shFE0A762E;
    weight_b_mem[ 608] = 32'shFB6C04B0;
    weight_b_mem[ 609] = 32'sh04625800;
    weight_b_mem[ 610] = 32'sh014CAA48;
    weight_b_mem[ 611] = 32'shFFC23390;
    weight_b_mem[ 612] = 32'sh04C53AE8;
    weight_b_mem[ 613] = 32'shFCAF9B64;
    weight_b_mem[ 614] = 32'shFAC619F8;
    weight_b_mem[ 615] = 32'shFF276F7A;
    weight_b_mem[ 616] = 32'shFF0280FD;
    weight_b_mem[ 617] = 32'sh03241FB4;
    weight_b_mem[ 618] = 32'shFE5BF3F6;
    weight_b_mem[ 619] = 32'shFB9A4D38;
    weight_b_mem[ 620] = 32'shFA7D3D18;
    weight_b_mem[ 621] = 32'sh0655F2F8;
    weight_b_mem[ 622] = 32'sh02E25D2C;
    weight_b_mem[ 623] = 32'shFC5F3E44;
    weight_b_mem[ 624] = 32'sh054A1648;
    weight_b_mem[ 625] = 32'shFFF8DC28;
    weight_b_mem[ 626] = 32'sh019A51CE;
    weight_b_mem[ 627] = 32'shFC94211C;
    weight_b_mem[ 628] = 32'shFAD753B0;
    weight_b_mem[ 629] = 32'shFD5E7090;
    weight_b_mem[ 630] = 32'shFCEE241C;
    weight_b_mem[ 631] = 32'sh02A26B90;
    weight_b_mem[ 632] = 32'sh0261A2E0;
    weight_b_mem[ 633] = 32'sh05A13B78;
    weight_b_mem[ 634] = 32'sh037831EC;
    weight_b_mem[ 635] = 32'shFC85E5EC;
    weight_b_mem[ 636] = 32'shF93C09E0;
    weight_b_mem[ 637] = 32'shFB54EB40;
    weight_b_mem[ 638] = 32'sh02BD42B0;
    weight_b_mem[ 639] = 32'sh00BA23F5;
    weight_b_mem[ 640] = 32'shFAFD0B38;
    weight_b_mem[ 641] = 32'sh01238DBA;
    weight_b_mem[ 642] = 32'sh05AB0E80;
    weight_b_mem[ 643] = 32'sh051A3F78;
    weight_b_mem[ 644] = 32'shFFD15FE2;
    weight_b_mem[ 645] = 32'sh0616A3C8;
    weight_b_mem[ 646] = 32'sh04D11A08;
    weight_b_mem[ 647] = 32'shFAA75D68;
    weight_b_mem[ 648] = 32'shFAD7CB10;
    weight_b_mem[ 649] = 32'shFA4717A8;
    weight_b_mem[ 650] = 32'sh03FBDE94;
    weight_b_mem[ 651] = 32'shFBB76258;
    weight_b_mem[ 652] = 32'sh00A59FEB;
    weight_b_mem[ 653] = 32'shFCA1DF48;
    weight_b_mem[ 654] = 32'sh045A65C0;
    weight_b_mem[ 655] = 32'sh00D95267;
    weight_b_mem[ 656] = 32'shFC1543DC;
    weight_b_mem[ 657] = 32'shFBF03278;
    weight_b_mem[ 658] = 32'sh05E71898;
    weight_b_mem[ 659] = 32'sh05A6D458;
    weight_b_mem[ 660] = 32'shFA9A6E70;
    weight_b_mem[ 661] = 32'sh036DE6B0;
    weight_b_mem[ 662] = 32'sh00564004;
    weight_b_mem[ 663] = 32'sh063DF5E0;
    weight_b_mem[ 664] = 32'shFFC343D6;
    weight_b_mem[ 665] = 32'sh07201120;
    weight_b_mem[ 666] = 32'shFC6E18DC;
    weight_b_mem[ 667] = 32'shFEC1FF32;
    weight_b_mem[ 668] = 32'shFF37D0A4;
    weight_b_mem[ 669] = 32'sh01AD570A;
    weight_b_mem[ 670] = 32'shFB013C10;
    weight_b_mem[ 671] = 32'sh032F49DC;
    weight_b_mem[ 672] = 32'shF8991BF0;
    weight_b_mem[ 673] = 32'shFE114DE8;
    weight_b_mem[ 674] = 32'sh0948AFE0;
    weight_b_mem[ 675] = 32'shFE97E0C8;
    weight_b_mem[ 676] = 32'shFD8CED34;
    weight_b_mem[ 677] = 32'sh01EBF812;
    weight_b_mem[ 678] = 32'sh01A5C3C2;
    weight_b_mem[ 679] = 32'shFF2EC284;
    weight_b_mem[ 680] = 32'shF7DF95A0;
    weight_b_mem[ 681] = 32'sh000ED2D0;
    weight_b_mem[ 682] = 32'sh01B9F986;
    weight_b_mem[ 683] = 32'sh01AE9CA0;
    weight_b_mem[ 684] = 32'sh0140E332;
    weight_b_mem[ 685] = 32'shFF86FA5A;
    weight_b_mem[ 686] = 32'shF9779D00;
    weight_b_mem[ 687] = 32'sh0879F9D0;
    weight_b_mem[ 688] = 32'sh019B519E;
    weight_b_mem[ 689] = 32'sh032AF55C;
    weight_b_mem[ 690] = 32'sh013E4344;
    weight_b_mem[ 691] = 32'shFCE84294;
    weight_b_mem[ 692] = 32'shFC332854;
    weight_b_mem[ 693] = 32'sh01552D3E;
    weight_b_mem[ 694] = 32'shFE93AF6E;
    weight_b_mem[ 695] = 32'sh06AFD2D0;
    weight_b_mem[ 696] = 32'shFFDD0CDD;
    weight_b_mem[ 697] = 32'shFBC9B748;
    weight_b_mem[ 698] = 32'shF8ACDC40;
    weight_b_mem[ 699] = 32'sh022688B0;
    weight_b_mem[ 700] = 32'sh043B56C0;
    weight_b_mem[ 701] = 32'shFC4955B4;
    weight_b_mem[ 702] = 32'shF87470E0;
    weight_b_mem[ 703] = 32'shFEFE89C8;
    weight_b_mem[ 704] = 32'sh0169D76C;
    weight_b_mem[ 705] = 32'sh027D29D8;
    weight_b_mem[ 706] = 32'shFE2E493E;
    weight_b_mem[ 707] = 32'shFEB7D1FE;
    weight_b_mem[ 708] = 32'sh02C311BC;
    weight_b_mem[ 709] = 32'shFD958E78;
    weight_b_mem[ 710] = 32'shFE43F432;
    weight_b_mem[ 711] = 32'sh057C12A0;
    weight_b_mem[ 712] = 32'shFBF15940;
    weight_b_mem[ 713] = 32'sh0184345C;
    weight_b_mem[ 714] = 32'shFE941682;
    weight_b_mem[ 715] = 32'sh035CA90C;
    weight_b_mem[ 716] = 32'sh03FF1F88;
    weight_b_mem[ 717] = 32'sh032CA6E0;
    weight_b_mem[ 718] = 32'sh05FB4EB8;
    weight_b_mem[ 719] = 32'sh002F6E8A;
    weight_b_mem[ 720] = 32'shF912CB78;
    weight_b_mem[ 721] = 32'shFD900D78;
    weight_b_mem[ 722] = 32'shFEFF0EC6;
    weight_b_mem[ 723] = 32'shFD0136E4;
    weight_b_mem[ 724] = 32'sh02CBB65C;
    weight_b_mem[ 725] = 32'shFFD4FC10;
    weight_b_mem[ 726] = 32'sh00915194;
    weight_b_mem[ 727] = 32'shFFAF79FD;
    weight_b_mem[ 728] = 32'sh01E450E4;
    weight_b_mem[ 729] = 32'shFACC5388;
    weight_b_mem[ 730] = 32'sh00BB075B;
    weight_b_mem[ 731] = 32'sh022241B0;
    weight_b_mem[ 732] = 32'shFCB242D0;
    weight_b_mem[ 733] = 32'sh01B035D4;
    weight_b_mem[ 734] = 32'shFBB2FFB0;
    weight_b_mem[ 735] = 32'shFAD83268;
    weight_b_mem[ 736] = 32'sh02E72438;
    weight_b_mem[ 737] = 32'sh014D4616;
    weight_b_mem[ 738] = 32'sh05DE0BD0;
    weight_b_mem[ 739] = 32'sh000204D2;
    weight_b_mem[ 740] = 32'sh002A194A;
    weight_b_mem[ 741] = 32'sh0708C770;
    weight_b_mem[ 742] = 32'sh07560810;
    weight_b_mem[ 743] = 32'sh05B8A2F0;
    weight_b_mem[ 744] = 32'shFD5F2850;
    weight_b_mem[ 745] = 32'sh00FFB317;
    weight_b_mem[ 746] = 32'sh06FB8D48;
    weight_b_mem[ 747] = 32'shFD37CBA4;
    weight_b_mem[ 748] = 32'sh0231139C;
    weight_b_mem[ 749] = 32'shFE62953E;
    weight_b_mem[ 750] = 32'shFA073DB0;
    weight_b_mem[ 751] = 32'sh056F78C0;
    weight_b_mem[ 752] = 32'shFB757828;
    weight_b_mem[ 753] = 32'sh059EA828;
    weight_b_mem[ 754] = 32'sh01C2F6AC;
    weight_b_mem[ 755] = 32'sh03DB17D4;
    weight_b_mem[ 756] = 32'sh0216F294;
    weight_b_mem[ 757] = 32'sh06C93DE0;
    weight_b_mem[ 758] = 32'shFBB6D600;
    weight_b_mem[ 759] = 32'sh01D5ECA6;
    weight_b_mem[ 760] = 32'shFBEF7F90;
    weight_b_mem[ 761] = 32'shFF5F8D8E;
    weight_b_mem[ 762] = 32'shFBAEC0B8;
    weight_b_mem[ 763] = 32'shFD749080;
    weight_b_mem[ 764] = 32'shFFC2DC80;
    weight_b_mem[ 765] = 32'sh00D11B83;
    weight_b_mem[ 766] = 32'sh04C631F0;
    weight_b_mem[ 767] = 32'shFF58E056;
    weight_b_mem[ 768] = 32'shFDBDAD90;
    weight_b_mem[ 769] = 32'sh0137F184;
    weight_b_mem[ 770] = 32'sh02354C44;
    weight_b_mem[ 771] = 32'shFF34EFB1;
    weight_b_mem[ 772] = 32'sh005E9ABB;
    weight_b_mem[ 773] = 32'shF96A8A18;
    weight_b_mem[ 774] = 32'sh0391D8B4;
    weight_b_mem[ 775] = 32'sh04FF4FA8;
    weight_b_mem[ 776] = 32'sh037A2BC8;
    weight_b_mem[ 777] = 32'sh033BB428;
    weight_b_mem[ 778] = 32'sh024F859C;
    weight_b_mem[ 779] = 32'shFDCE37F0;
    weight_b_mem[ 780] = 32'sh0245D6C4;
    weight_b_mem[ 781] = 32'sh01D0DA3E;
    weight_b_mem[ 782] = 32'sh05844AE0;
    weight_b_mem[ 783] = 32'shFDDC8F1C;
    weight_b_mem[ 784] = 32'shFE0AEC52;
    weight_b_mem[ 785] = 32'sh008A089F;
    weight_b_mem[ 786] = 32'sh0197D96E;
    weight_b_mem[ 787] = 32'shFD506D48;
    weight_b_mem[ 788] = 32'shFF2BEB08;
    weight_b_mem[ 789] = 32'sh07C40DD0;
    weight_b_mem[ 790] = 32'shFDCBA8C8;
    weight_b_mem[ 791] = 32'shFDAE7F88;
    weight_b_mem[ 792] = 32'shFEE0A33A;
    weight_b_mem[ 793] = 32'shFA7741A8;
    weight_b_mem[ 794] = 32'shFD05B5A0;
    weight_b_mem[ 795] = 32'sh053DBBA8;
    weight_b_mem[ 796] = 32'sh000D2836;
    weight_b_mem[ 797] = 32'sh0132DC20;
    weight_b_mem[ 798] = 32'sh0376C2DC;
    weight_b_mem[ 799] = 32'sh08289920;
    weight_b_mem[ 800] = 32'sh02658A4C;
    weight_b_mem[ 801] = 32'sh04B7FF70;
    weight_b_mem[ 802] = 32'sh07DAE970;
    weight_b_mem[ 803] = 32'sh0160A976;
    weight_b_mem[ 804] = 32'sh0574F7A0;
    weight_b_mem[ 805] = 32'shFF85306D;
    weight_b_mem[ 806] = 32'shFE5FFF4C;
    weight_b_mem[ 807] = 32'shFBDBB890;
    weight_b_mem[ 808] = 32'shFF95EBC3;
    weight_b_mem[ 809] = 32'sh02C67F88;
    weight_b_mem[ 810] = 32'shFC56F2B0;
    weight_b_mem[ 811] = 32'sh06F7C108;
    weight_b_mem[ 812] = 32'shFC39598C;
    weight_b_mem[ 813] = 32'shFC7009C0;
    weight_b_mem[ 814] = 32'shFCC9A5E0;
    weight_b_mem[ 815] = 32'shFF08B926;
    weight_b_mem[ 816] = 32'sh020C754C;
    weight_b_mem[ 817] = 32'shFAB3A550;
    weight_b_mem[ 818] = 32'shFF4E4F52;
    weight_b_mem[ 819] = 32'sh035DBA5C;
    weight_b_mem[ 820] = 32'shFDAAE558;
    weight_b_mem[ 821] = 32'sh00B7BF2B;
    weight_b_mem[ 822] = 32'shFE8D7760;
    weight_b_mem[ 823] = 32'sh01770BE6;
    weight_b_mem[ 824] = 32'sh00EF5310;
    weight_b_mem[ 825] = 32'sh04917FA0;
    weight_b_mem[ 826] = 32'shF9D50838;
    weight_b_mem[ 827] = 32'shFD853F3C;
    weight_b_mem[ 828] = 32'sh02F7C828;
    weight_b_mem[ 829] = 32'sh06633C00;
    weight_b_mem[ 830] = 32'shFED739BA;
    weight_b_mem[ 831] = 32'sh04471E70;
    weight_b_mem[ 832] = 32'shFED951E0;
    weight_b_mem[ 833] = 32'sh034B4A50;
    weight_b_mem[ 834] = 32'shFD6A3BC0;
    weight_b_mem[ 835] = 32'shFF87E984;
    weight_b_mem[ 836] = 32'sh03E1CB74;
    weight_b_mem[ 837] = 32'sh0286FAFC;
    weight_b_mem[ 838] = 32'sh0CB627D0;
    weight_b_mem[ 839] = 32'sh03AD20B0;
    weight_b_mem[ 840] = 32'sh006709A8;
    weight_b_mem[ 841] = 32'sh012DDA8A;
    weight_b_mem[ 842] = 32'sh01329B02;
    weight_b_mem[ 843] = 32'sh0BD6FB40;
    weight_b_mem[ 844] = 32'shFDA1551C;
    weight_b_mem[ 845] = 32'sh001B0855;
    weight_b_mem[ 846] = 32'shFC98199C;
    weight_b_mem[ 847] = 32'sh04245D28;
    weight_b_mem[ 848] = 32'sh01CC13A4;
    weight_b_mem[ 849] = 32'sh02F2DA34;
    weight_b_mem[ 850] = 32'shF9BED3D0;
    weight_b_mem[ 851] = 32'sh0075B183;
    weight_b_mem[ 852] = 32'sh0A2208B0;
    weight_b_mem[ 853] = 32'sh0B4EB3B0;
    weight_b_mem[ 854] = 32'sh0ADEBA90;
    weight_b_mem[ 855] = 32'shFE67FA26;
    weight_b_mem[ 856] = 32'sh0DE34A70;
    weight_b_mem[ 857] = 32'shF6BBEA70;
    weight_b_mem[ 858] = 32'shFB7B3C10;
    weight_b_mem[ 859] = 32'sh08F43E20;
    weight_b_mem[ 860] = 32'shFE2F4B94;
    weight_b_mem[ 861] = 32'sh03F1FCEC;
    weight_b_mem[ 862] = 32'sh02D77754;
    weight_b_mem[ 863] = 32'sh0399CBA8;
    weight_b_mem[ 864] = 32'sh01726D26;
    weight_b_mem[ 865] = 32'sh029C0C2C;
    weight_b_mem[ 866] = 32'shF8B10D48;
    weight_b_mem[ 867] = 32'sh01CE5872;
    weight_b_mem[ 868] = 32'sh04D2E320;
    weight_b_mem[ 869] = 32'sh06900D18;
    weight_b_mem[ 870] = 32'sh020E07F8;
    weight_b_mem[ 871] = 32'shFEEA7E52;
    weight_b_mem[ 872] = 32'shFE44A572;
    weight_b_mem[ 873] = 32'shFF394556;
    weight_b_mem[ 874] = 32'shFE30D57C;
    weight_b_mem[ 875] = 32'shFB511DA0;
    weight_b_mem[ 876] = 32'sh02F640E8;
    weight_b_mem[ 877] = 32'shFED88F5C;
    weight_b_mem[ 878] = 32'shFC77F90C;
    weight_b_mem[ 879] = 32'sh08380A20;
    weight_b_mem[ 880] = 32'sh03A0F42C;
    weight_b_mem[ 881] = 32'shF7411510;
    weight_b_mem[ 882] = 32'sh0988D0F0;
    weight_b_mem[ 883] = 32'sh02A048EC;
    weight_b_mem[ 884] = 32'sh005A8C4A;
    weight_b_mem[ 885] = 32'shFE70DBD0;
    weight_b_mem[ 886] = 32'shFE4445F8;
    weight_b_mem[ 887] = 32'shFFEA7A23;
    weight_b_mem[ 888] = 32'shEA675A60;
    weight_b_mem[ 889] = 32'sh08213A60;
    weight_b_mem[ 890] = 32'shFD367488;
    weight_b_mem[ 891] = 32'shF9A479F0;
    weight_b_mem[ 892] = 32'shFB0759B0;
    weight_b_mem[ 893] = 32'sh05ADC140;
    weight_b_mem[ 894] = 32'sh05A5F130;
    weight_b_mem[ 895] = 32'sh00385415;
    weight_b_mem[ 896] = 32'shF9137520;
    weight_b_mem[ 897] = 32'shFC817938;
    weight_b_mem[ 898] = 32'shFCCA6D4C;
    weight_b_mem[ 899] = 32'sh00F23390;
    weight_b_mem[ 900] = 32'shFC5003C8;
    weight_b_mem[ 901] = 32'sh03FC10F0;
    weight_b_mem[ 902] = 32'shF6035F30;
    weight_b_mem[ 903] = 32'sh001409D3;
    weight_b_mem[ 904] = 32'shFBCDC468;
    weight_b_mem[ 905] = 32'shFD6D5CC8;
    weight_b_mem[ 906] = 32'sh04B7C380;
    weight_b_mem[ 907] = 32'sh0607E978;
    weight_b_mem[ 908] = 32'sh028A1830;
    weight_b_mem[ 909] = 32'sh013D9420;
    weight_b_mem[ 910] = 32'shFA2A2940;
    weight_b_mem[ 911] = 32'shFFABDE2A;
    weight_b_mem[ 912] = 32'shFD16E158;
    weight_b_mem[ 913] = 32'shFECDBEE0;
    weight_b_mem[ 914] = 32'sh03A3CDBC;
    weight_b_mem[ 915] = 32'sh042FFE78;
    weight_b_mem[ 916] = 32'shFDF00D4C;
    weight_b_mem[ 917] = 32'shFBA00E98;
    weight_b_mem[ 918] = 32'sh0B49EAE0;
    weight_b_mem[ 919] = 32'shFEE6BE7C;
    weight_b_mem[ 920] = 32'shFD2AAE30;
    weight_b_mem[ 921] = 32'sh0A70B620;
    weight_b_mem[ 922] = 32'shFE649CFC;
    weight_b_mem[ 923] = 32'shF5AC6A30;
    weight_b_mem[ 924] = 32'shFBE77E08;
    weight_b_mem[ 925] = 32'shFE2A6D1C;
    weight_b_mem[ 926] = 32'sh06508508;
    weight_b_mem[ 927] = 32'shFEA35854;
    weight_b_mem[ 928] = 32'sh0423D160;
    weight_b_mem[ 929] = 32'sh05512CF8;
    weight_b_mem[ 930] = 32'shFDCC777C;
    weight_b_mem[ 931] = 32'sh02AED8B0;
    weight_b_mem[ 932] = 32'sh0179E27E;
    weight_b_mem[ 933] = 32'shFEB721F6;
    weight_b_mem[ 934] = 32'shF9C1A830;
    weight_b_mem[ 935] = 32'shFED16DE8;
    weight_b_mem[ 936] = 32'sh04E0A290;
    weight_b_mem[ 937] = 32'shFB56F910;
    weight_b_mem[ 938] = 32'shFC3B8650;
    weight_b_mem[ 939] = 32'shFEBE2032;
    weight_b_mem[ 940] = 32'shFE2C398C;
    weight_b_mem[ 941] = 32'sh02AD0E04;
    weight_b_mem[ 942] = 32'sh01700DEC;
    weight_b_mem[ 943] = 32'shFFE6051E;
    weight_b_mem[ 944] = 32'sh00199D5C;
    weight_b_mem[ 945] = 32'shFEC7C066;
    weight_b_mem[ 946] = 32'shFEE42C78;
    weight_b_mem[ 947] = 32'sh01FC0944;
    weight_b_mem[ 948] = 32'sh04CC0F30;
    weight_b_mem[ 949] = 32'shFAFFE8A0;
    weight_b_mem[ 950] = 32'sh01EE8598;
    weight_b_mem[ 951] = 32'sh0297A7F4;
    weight_b_mem[ 952] = 32'sh08677300;
    weight_b_mem[ 953] = 32'shFBE31CD0;
    weight_b_mem[ 954] = 32'sh04C8DF88;
    weight_b_mem[ 955] = 32'shFDA0E7AC;
    weight_b_mem[ 956] = 32'sh02194AF0;
    weight_b_mem[ 957] = 32'shFF4B68FE;
    weight_b_mem[ 958] = 32'sh0755ADE8;
    weight_b_mem[ 959] = 32'sh00F642C4;
    weight_b_mem[ 960] = 32'shFD599158;
    weight_b_mem[ 961] = 32'shFEB99200;
    weight_b_mem[ 962] = 32'sh016C0DE0;
    weight_b_mem[ 963] = 32'shFB8F9828;
    weight_b_mem[ 964] = 32'shFF291233;
    weight_b_mem[ 965] = 32'sh00F68C32;
    weight_b_mem[ 966] = 32'shFB42AE08;
    weight_b_mem[ 967] = 32'shF93D1720;
    weight_b_mem[ 968] = 32'shFCD1F568;
    weight_b_mem[ 969] = 32'sh004567AA;
    weight_b_mem[ 970] = 32'sh040116A8;
    weight_b_mem[ 971] = 32'shFD071190;
    weight_b_mem[ 972] = 32'sh0099A0ED;
    weight_b_mem[ 973] = 32'shFFA9543E;
    weight_b_mem[ 974] = 32'sh023DD8E0;
    weight_b_mem[ 975] = 32'sh0163CFC8;
    weight_b_mem[ 976] = 32'shFFEBBF04;
    weight_b_mem[ 977] = 32'sh07ADA108;
    weight_b_mem[ 978] = 32'sh037A7C18;
    weight_b_mem[ 979] = 32'sh03D9F0F0;
    weight_b_mem[ 980] = 32'sh03438748;
    weight_b_mem[ 981] = 32'shF678A160;
    weight_b_mem[ 982] = 32'shFFF0894E;
    weight_b_mem[ 983] = 32'sh01F82FB4;
    weight_b_mem[ 984] = 32'sh054EE540;
    weight_b_mem[ 985] = 32'shEF9EAAC0;
    weight_b_mem[ 986] = 32'shFCBE00C0;
    weight_b_mem[ 987] = 32'sh09737060;
    weight_b_mem[ 988] = 32'sh030733AC;
    weight_b_mem[ 989] = 32'shFDF78EE8;
    weight_b_mem[ 990] = 32'sh0001468F;
    weight_b_mem[ 991] = 32'sh05889708;
    weight_b_mem[ 992] = 32'shFA8F0568;
    weight_b_mem[ 993] = 32'shFDF4C224;
    weight_b_mem[ 994] = 32'shFC5BDAA4;
    weight_b_mem[ 995] = 32'sh06169E78;
    weight_b_mem[ 996] = 32'sh017B401C;
    weight_b_mem[ 997] = 32'sh08395500;
    weight_b_mem[ 998] = 32'sh01B16F9C;
    weight_b_mem[ 999] = 32'sh04966B40;
    weight_b_mem[1000] = 32'shFDD713D8;
    weight_b_mem[1001] = 32'sh03AE8E0C;
    weight_b_mem[1002] = 32'sh0279F46C;
    weight_b_mem[1003] = 32'sh017520B4;
    weight_b_mem[1004] = 32'shFF0CF17B;
    weight_b_mem[1005] = 32'sh04010DE8;
    weight_b_mem[1006] = 32'shFF1FDDAD;
    weight_b_mem[1007] = 32'sh07579BE8;
    weight_b_mem[1008] = 32'shFE487F08;
    weight_b_mem[1009] = 32'shFC118BE8;
    weight_b_mem[1010] = 32'sh00C333F9;
    weight_b_mem[1011] = 32'shFF23895B;
    weight_b_mem[1012] = 32'shFEB5F540;
    weight_b_mem[1013] = 32'sh011819F2;
    weight_b_mem[1014] = 32'sh06331C08;
    weight_b_mem[1015] = 32'shFED9C84C;
    weight_b_mem[1016] = 32'sh06F0A168;
    weight_b_mem[1017] = 32'shFB171B08;
    weight_b_mem[1018] = 32'sh004ACD3E;
    weight_b_mem[1019] = 32'sh03712244;
    weight_b_mem[1020] = 32'shFDDBA9CC;
    weight_b_mem[1021] = 32'sh0348BDA4;
    weight_b_mem[1022] = 32'shFC9CC134;
    weight_b_mem[1023] = 32'shFD75AEB0;
    weight_b_mem[1024] = 32'shFC895A6C;
    weight_b_mem[1025] = 32'sh005536E3;
    weight_b_mem[1026] = 32'sh034B0D00;
    weight_b_mem[1027] = 32'sh017B5CA8;
    weight_b_mem[1028] = 32'sh02FC5564;
    weight_b_mem[1029] = 32'sh0281D544;
    weight_b_mem[1030] = 32'sh02F5A8B8;
    weight_b_mem[1031] = 32'shFC2F675C;
    weight_b_mem[1032] = 32'shFF5B5187;
    weight_b_mem[1033] = 32'shFA73A060;
    weight_b_mem[1034] = 32'shFED1F91C;
    weight_b_mem[1035] = 32'shFD5FE500;
    weight_b_mem[1036] = 32'shFD61E3AC;
    weight_b_mem[1037] = 32'shFC473CD0;
    weight_b_mem[1038] = 32'sh0322CA98;
    weight_b_mem[1039] = 32'sh02173FB0;
    weight_b_mem[1040] = 32'sh0507A2D0;
    weight_b_mem[1041] = 32'sh01B22E3A;
    weight_b_mem[1042] = 32'sh01DFE6CE;
    weight_b_mem[1043] = 32'sh059E03A0;
    weight_b_mem[1044] = 32'sh0186E2AA;
    weight_b_mem[1045] = 32'sh03C316E0;
    weight_b_mem[1046] = 32'sh03304A64;
    weight_b_mem[1047] = 32'shFE8804B8;
    weight_b_mem[1048] = 32'shFEED3C32;
    weight_b_mem[1049] = 32'shFED85300;
    weight_b_mem[1050] = 32'shFAA72C30;
    weight_b_mem[1051] = 32'shFEB5E90A;
    weight_b_mem[1052] = 32'shFE52B66C;
    weight_b_mem[1053] = 32'sh028701B0;
    weight_b_mem[1054] = 32'sh00E2A2E1;
    weight_b_mem[1055] = 32'sh000BF0C5;
    weight_b_mem[1056] = 32'sh0942CCE0;
    weight_b_mem[1057] = 32'shFF157B1A;
    weight_b_mem[1058] = 32'sh059A4968;
    weight_b_mem[1059] = 32'sh0163A80A;
    weight_b_mem[1060] = 32'shFCE0A540;
    weight_b_mem[1061] = 32'shFD0F1FE0;
    weight_b_mem[1062] = 32'sh088C08B0;
    weight_b_mem[1063] = 32'shFF86D2CF;
    weight_b_mem[1064] = 32'shFDE02CA8;
    weight_b_mem[1065] = 32'sh018C64E0;
    weight_b_mem[1066] = 32'sh01C93D18;
    weight_b_mem[1067] = 32'shFE7477BC;
    weight_b_mem[1068] = 32'sh066A6BD8;
    weight_b_mem[1069] = 32'shFDF7FE94;
    weight_b_mem[1070] = 32'sh002E53FC;
    weight_b_mem[1071] = 32'sh06D71328;
    weight_b_mem[1072] = 32'shFED2CA48;
    weight_b_mem[1073] = 32'sh041A6040;
    weight_b_mem[1074] = 32'sh050062E8;
    weight_b_mem[1075] = 32'shFF454A51;
    weight_b_mem[1076] = 32'shF88E4E08;
    weight_b_mem[1077] = 32'shFF45A1D5;
    weight_b_mem[1078] = 32'sh06C2A118;
    weight_b_mem[1079] = 32'shFFAA4B90;
    weight_b_mem[1080] = 32'shFB1FDFC0;
    weight_b_mem[1081] = 32'sh025CE7E0;
    weight_b_mem[1082] = 32'shFAB3C4F8;
    weight_b_mem[1083] = 32'shFB315FB0;
    weight_b_mem[1084] = 32'sh059193C8;
    weight_b_mem[1085] = 32'shFB592638;
    weight_b_mem[1086] = 32'shFD8B6EA8;
    weight_b_mem[1087] = 32'shFFD5C079;
    weight_b_mem[1088] = 32'shFEDC0E58;
    weight_b_mem[1089] = 32'sh033D9F04;
    weight_b_mem[1090] = 32'shFFAAB7F2;
    weight_b_mem[1091] = 32'shFE786B28;
    weight_b_mem[1092] = 32'sh02824020;
    weight_b_mem[1093] = 32'sh0835B500;
    weight_b_mem[1094] = 32'sh0808F020;
    weight_b_mem[1095] = 32'sh03BC17F8;
    weight_b_mem[1096] = 32'sh0739F5C8;
    weight_b_mem[1097] = 32'sh03626C68;
    weight_b_mem[1098] = 32'shFE944C8E;
    weight_b_mem[1099] = 32'shFA616AB8;
    weight_b_mem[1100] = 32'shFF3B9871;
    weight_b_mem[1101] = 32'shFDD05C04;
    weight_b_mem[1102] = 32'sh06CB0D58;
    weight_b_mem[1103] = 32'shFAC39F28;
    weight_b_mem[1104] = 32'sh00AC015C;
    weight_b_mem[1105] = 32'sh0160047E;
    weight_b_mem[1106] = 32'sh056476A8;
    weight_b_mem[1107] = 32'sh009727E6;
    weight_b_mem[1108] = 32'shF9FB8AF0;
    weight_b_mem[1109] = 32'shFB087EE0;
    weight_b_mem[1110] = 32'sh037AE69C;
    weight_b_mem[1111] = 32'sh02F5A008;
    weight_b_mem[1112] = 32'shFECD7ADE;
    weight_b_mem[1113] = 32'shFD3E3B30;
    weight_b_mem[1114] = 32'sh03707AA8;
    weight_b_mem[1115] = 32'shFD63B474;
    weight_b_mem[1116] = 32'shFABA0528;
    weight_b_mem[1117] = 32'shFD951AD0;
    weight_b_mem[1118] = 32'shFF68BCCC;
    weight_b_mem[1119] = 32'shF89934F8;
    weight_b_mem[1120] = 32'shFB3AB588;
    weight_b_mem[1121] = 32'sh001AA26E;
    weight_b_mem[1122] = 32'shFA3C6C40;
    weight_b_mem[1123] = 32'shFF26BF5C;
    weight_b_mem[1124] = 32'shFE0843B6;
    weight_b_mem[1125] = 32'sh04ECF2F8;
    weight_b_mem[1126] = 32'shF90ABE98;
    weight_b_mem[1127] = 32'shFB705FF8;
    weight_b_mem[1128] = 32'shFEFE0F7A;
    weight_b_mem[1129] = 32'sh05BFC600;
    weight_b_mem[1130] = 32'sh059DFCE0;
    weight_b_mem[1131] = 32'sh086F3C50;
    weight_b_mem[1132] = 32'sh0225F744;
    weight_b_mem[1133] = 32'sh0725C908;
    weight_b_mem[1134] = 32'shFE31364E;
    weight_b_mem[1135] = 32'sh05485250;
    weight_b_mem[1136] = 32'shFA474DF0;
    weight_b_mem[1137] = 32'shFA2E6900;
    weight_b_mem[1138] = 32'sh06A32A90;
    weight_b_mem[1139] = 32'sh06478C98;
    weight_b_mem[1140] = 32'sh06CB67C0;
    weight_b_mem[1141] = 32'shFB105D40;
    weight_b_mem[1142] = 32'shFEA88374;
    weight_b_mem[1143] = 32'shFF86D8BB;
    weight_b_mem[1144] = 32'shFDDA3478;
    weight_b_mem[1145] = 32'sh05BC5458;
    weight_b_mem[1146] = 32'sh00858AD4;
    weight_b_mem[1147] = 32'sh081D6180;
    weight_b_mem[1148] = 32'shFA63CAC0;
    weight_b_mem[1149] = 32'sh007E419C;
    weight_b_mem[1150] = 32'shF9C49058;
    weight_b_mem[1151] = 32'sh00935687;
    weight_b_mem[1152] = 32'shFE3FC3CC;
    weight_b_mem[1153] = 32'shFD83A70C;
    weight_b_mem[1154] = 32'shFFC326E5;
    weight_b_mem[1155] = 32'sh010BC00C;
    weight_b_mem[1156] = 32'shFFE8EEA4;
    weight_b_mem[1157] = 32'sh0144C4B8;
    weight_b_mem[1158] = 32'shFE7D2382;
    weight_b_mem[1159] = 32'shFE7FB7B4;
    weight_b_mem[1160] = 32'shFDD57984;
    weight_b_mem[1161] = 32'shFF953952;
    weight_b_mem[1162] = 32'shFFDBE8C1;
    weight_b_mem[1163] = 32'shFD053E04;
    weight_b_mem[1164] = 32'sh015CE2CE;
    weight_b_mem[1165] = 32'shFD7B8788;
    weight_b_mem[1166] = 32'sh0398B7E0;
    weight_b_mem[1167] = 32'shFEA97BE6;
    weight_b_mem[1168] = 32'sh00C952D1;
    weight_b_mem[1169] = 32'shFDA0AD60;
    weight_b_mem[1170] = 32'shFEC741E4;
    weight_b_mem[1171] = 32'shFF460980;
    weight_b_mem[1172] = 32'sh0038E453;
    weight_b_mem[1173] = 32'shFF53E6F8;
    weight_b_mem[1174] = 32'sh011D421E;
    weight_b_mem[1175] = 32'sh010FED18;
    weight_b_mem[1176] = 32'sh0194F34C;
    weight_b_mem[1177] = 32'sh02F2BBB8;
    weight_b_mem[1178] = 32'shFD355514;
    weight_b_mem[1179] = 32'shFDEC2F9C;
    weight_b_mem[1180] = 32'shFC974B4C;
    weight_b_mem[1181] = 32'shFE363EA6;
    weight_b_mem[1182] = 32'shFF995DAA;
    weight_b_mem[1183] = 32'sh021D0CC0;
    weight_b_mem[1184] = 32'sh042B3BC8;
    weight_b_mem[1185] = 32'sh02AC1F28;
    weight_b_mem[1186] = 32'shF9803368;
    weight_b_mem[1187] = 32'shFBACB3E8;
    weight_b_mem[1188] = 32'sh04F010D0;
    weight_b_mem[1189] = 32'shFDF61324;
    weight_b_mem[1190] = 32'shFEDD27D2;
    weight_b_mem[1191] = 32'shFAC5F290;
    weight_b_mem[1192] = 32'sh02BF0AE4;
    weight_b_mem[1193] = 32'sh0A64E8A0;
    weight_b_mem[1194] = 32'shFC5C8A8C;
    weight_b_mem[1195] = 32'sh0477C908;
    weight_b_mem[1196] = 32'sh09BB57C0;
    weight_b_mem[1197] = 32'sh058D6FB0;
    weight_b_mem[1198] = 32'shF872A768;
    weight_b_mem[1199] = 32'sh05CB5A78;
    weight_b_mem[1200] = 32'sh05125D18;
    weight_b_mem[1201] = 32'sh03556C4C;
    weight_b_mem[1202] = 32'sh04014A58;
    weight_b_mem[1203] = 32'sh0704DF38;
    weight_b_mem[1204] = 32'shFD0C44CC;
    weight_b_mem[1205] = 32'sh017E82FA;
    weight_b_mem[1206] = 32'shFC535760;
    weight_b_mem[1207] = 32'shF84D1728;
    weight_b_mem[1208] = 32'shFAE58808;
    weight_b_mem[1209] = 32'shFCC4A580;
    weight_b_mem[1210] = 32'shF8AC50D8;
    weight_b_mem[1211] = 32'shFE54F202;
    weight_b_mem[1212] = 32'sh00955726;
    weight_b_mem[1213] = 32'sh053EF2D0;
    weight_b_mem[1214] = 32'sh038CC4C4;
    weight_b_mem[1215] = 32'shFEC1A3CC;
    weight_b_mem[1216] = 32'shF987C6C8;
    weight_b_mem[1217] = 32'shF9F70F18;
    weight_b_mem[1218] = 32'shFE117B14;
    weight_b_mem[1219] = 32'shFB8F2A38;
    weight_b_mem[1220] = 32'shFCAFC718;
    weight_b_mem[1221] = 32'shFD40349C;
    weight_b_mem[1222] = 32'shFD4E3E08;
    weight_b_mem[1223] = 32'sh031EDB00;
    weight_b_mem[1224] = 32'shFCA77874;
    weight_b_mem[1225] = 32'sh0379D2B0;
    weight_b_mem[1226] = 32'shFAC2BEB8;
    weight_b_mem[1227] = 32'sh0246F950;
    weight_b_mem[1228] = 32'shFE7C05D0;
    weight_b_mem[1229] = 32'sh03389778;
    weight_b_mem[1230] = 32'shFF2D2A85;
    weight_b_mem[1231] = 32'sh044BFCB0;
    weight_b_mem[1232] = 32'sh011E9B40;
    weight_b_mem[1233] = 32'sh035DAD30;
    weight_b_mem[1234] = 32'sh05BD8358;
    weight_b_mem[1235] = 32'sh033EFD1C;
    weight_b_mem[1236] = 32'sh060B4410;
    weight_b_mem[1237] = 32'sh00F9799A;
    weight_b_mem[1238] = 32'shFC84FB8C;
    weight_b_mem[1239] = 32'sh013D8982;
    weight_b_mem[1240] = 32'sh0484BF38;
    weight_b_mem[1241] = 32'shFCB224D0;
    weight_b_mem[1242] = 32'sh031C787C;
    weight_b_mem[1243] = 32'sh04A35450;
    weight_b_mem[1244] = 32'shF9B9B358;
    weight_b_mem[1245] = 32'sh025BBC4C;
    weight_b_mem[1246] = 32'sh02A93530;
    weight_b_mem[1247] = 32'shFD3ABF1C;
    weight_b_mem[1248] = 32'shFC279DC8;
    weight_b_mem[1249] = 32'sh04B082C8;
    weight_b_mem[1250] = 32'sh05E12E88;
    weight_b_mem[1251] = 32'shFF9D9EC8;
    weight_b_mem[1252] = 32'shFF836CFC;
    weight_b_mem[1253] = 32'shFEC70EE0;
    weight_b_mem[1254] = 32'sh0446FD58;
    weight_b_mem[1255] = 32'shFB13B8F8;
    weight_b_mem[1256] = 32'shFB49A160;
    weight_b_mem[1257] = 32'shFDABB8A0;
    weight_b_mem[1258] = 32'shFFC2577E;
    weight_b_mem[1259] = 32'sh04AE7A60;
    weight_b_mem[1260] = 32'shF9EF3E10;
    weight_b_mem[1261] = 32'sh00CA798D;
    weight_b_mem[1262] = 32'sh03503D6C;
    weight_b_mem[1263] = 32'shFE66CA04;
    weight_b_mem[1264] = 32'sh02FED0E4;
    weight_b_mem[1265] = 32'sh04AC1178;
    weight_b_mem[1266] = 32'sh05EF7CA0;
    weight_b_mem[1267] = 32'shFBF8AB88;
    weight_b_mem[1268] = 32'sh023727AC;
    weight_b_mem[1269] = 32'sh074D5248;
    weight_b_mem[1270] = 32'sh05B51990;
    weight_b_mem[1271] = 32'sh0404F0A0;
    weight_b_mem[1272] = 32'sh02A63800;
    weight_b_mem[1273] = 32'sh0366B7EC;
    weight_b_mem[1274] = 32'sh06CD8318;
    weight_b_mem[1275] = 32'sh041FBB00;
    weight_b_mem[1276] = 32'shFF6632A6;
    weight_b_mem[1277] = 32'shFC85CFFC;
    weight_b_mem[1278] = 32'shFF0D34DB;
    weight_b_mem[1279] = 32'sh04069D28;
    weight_b_mem[1280] = 32'shFF6EE13F;
    weight_b_mem[1281] = 32'sh0019E12D;
    weight_b_mem[1282] = 32'shFBE36CB0;
end
