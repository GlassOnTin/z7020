// sine_lut.v — Quarter-wave sine lookup table for SIREN activation
//
// Computes sin(angle) for Q4.28 fixed-point inputs and outputs.
// Uses 256-entry quarter-wave table with quadrant reconstruction.
//
// Input:  angle in Q4.28 radians (any value, reduced mod 2*pi)
// Output: sin(angle) in Q4.28 (range [-1, +1])
//
// Latency: 2 cycles (registered input + registered output)
//
// For SIREN networks, the activation is sin(omega * x) where omega
// is typically 30.0 for the first layer and 1.0 for hidden layers.
// The omega scaling is done in the MLP core before calling this LUT.

`timescale 1ns / 1ps

module sine_lut #(
    parameter WIDTH = 32,
    parameter FRAC  = 28
)(
    input  wire                    clk,
    input  wire signed [WIDTH-1:0] angle,   // Q4.28 radians
    output reg  signed [WIDTH-1:0] result   // Q4.28 sin(angle)
);

    // =========================================================
    // Constants in Q4.28
    // =========================================================
    // pi   = 3.14159265... * 2^28 = 843314857  = 32'h3243_F6A9
    // 2*pi = 6.28318530... * 2^28 = 1686629713 = 32'h6487_ED51
    // pi/2 = 1.57079632... * 2^28 = 421657428  = 32'h1921_FB54
    localparam signed [WIDTH-1:0] TWO_PI  = 32'sh6487_ED51;
    localparam signed [WIDTH-1:0] PI      = 32'sh3243_F6A9;
    localparam signed [WIDTH-1:0] HALF_PI = 32'sh1921_FB54;

    // =========================================================
    // Quarter-wave sine table: 256 entries for [0, pi/2)
    // =========================================================
    // Entry k = sin(k * pi/2 / 256) in Q4.28
    // sin(0) = 0, sin(pi/2) = 1.0 = 0x10000000
    //
    // Generated by: round(sin(k * pi / 512) * 2^28) for k=0..255
    reg signed [WIDTH-1:0] sine_table [0:255];

    // Table values: round(sin(k * pi / 512) * 2^28) for k=0..255
    // Range: [0, 0x0FFFEC43] representing [0.0, 0.99998] in Q4.28
    initial begin
        sine_table[  0] = 32'sh00000000; sine_table[  1] = 32'sh001921F1;
        sine_table[  2] = 32'sh003243A4; sine_table[  3] = 32'sh004B64DB;
        sine_table[  4] = 32'sh00648558; sine_table[  5] = 32'sh007DA4DD;
        sine_table[  6] = 32'sh0096C32C; sine_table[  7] = 32'sh00AFE007;
        sine_table[  8] = 32'sh00C8FB30; sine_table[  9] = 32'sh00E21469;
        sine_table[ 10] = 32'sh00FB2B74; sine_table[ 11] = 32'sh01144013;
        sine_table[ 12] = 32'sh012D5209; sine_table[ 13] = 32'sh01466118;
        sine_table[ 14] = 32'sh015F6D01; sine_table[ 15] = 32'sh01787587;
        sine_table[ 16] = 32'sh01917A6C; sine_table[ 17] = 32'sh01AA7B72;
        sine_table[ 18] = 32'sh01C3785C; sine_table[ 19] = 32'sh01DC70ED;
        sine_table[ 20] = 32'sh01F564E5; sine_table[ 21] = 32'sh020E5409;
        sine_table[ 22] = 32'sh02273E1A; sine_table[ 23] = 32'sh024022DB;
        sine_table[ 24] = 32'sh0259020E; sine_table[ 25] = 32'sh0271DB76;
        sine_table[ 26] = 32'sh028AAED6; sine_table[ 27] = 32'sh02A37BF1;
        sine_table[ 28] = 32'sh02BC4289; sine_table[ 29] = 32'sh02D50261;
        sine_table[ 30] = 32'sh02EDBB3C; sine_table[ 31] = 32'sh03066CDD;
        sine_table[ 32] = 32'sh031F1708; sine_table[ 33] = 32'sh0337B97E;
        sine_table[ 34] = 32'sh03505405; sine_table[ 35] = 32'sh0368E65E;
        sine_table[ 36] = 32'sh0381704D; sine_table[ 37] = 32'sh0399F196;
        sine_table[ 38] = 32'sh03B269FD; sine_table[ 39] = 32'sh03CAD944;
        sine_table[ 40] = 32'sh03E33F2F; sine_table[ 41] = 32'sh03FB9B83;
        sine_table[ 42] = 32'sh0413EE04; sine_table[ 43] = 32'sh042C3674;
        sine_table[ 44] = 32'sh04447499; sine_table[ 45] = 32'sh045CA836;
        sine_table[ 46] = 32'sh0474D110; sine_table[ 47] = 32'sh048CEEEB;
        sine_table[ 48] = 32'sh04A5018C; sine_table[ 49] = 32'sh04BD08B7;
        sine_table[ 50] = 32'sh04D50431; sine_table[ 51] = 32'sh04ECF3BF;
        sine_table[ 52] = 32'sh0504D725; sine_table[ 53] = 32'sh051CAE29;
        sine_table[ 54] = 32'sh05347891; sine_table[ 55] = 32'sh054C3620;
        sine_table[ 56] = 32'sh0563E69D; sine_table[ 57] = 32'sh057B89CE;
        sine_table[ 58] = 32'sh05931F77; sine_table[ 59] = 32'sh05AAA75F;
        sine_table[ 60] = 32'sh05C2214C; sine_table[ 61] = 32'sh05D98D04;
        sine_table[ 62] = 32'sh05F0EA4C; sine_table[ 63] = 32'sh060838EC;
        sine_table[ 64] = 32'sh061F78AA; sine_table[ 65] = 32'sh0636A94C;
        sine_table[ 66] = 32'sh064DCA99; sine_table[ 67] = 32'sh0664DC58;
        sine_table[ 68] = 32'sh067BDE51; sine_table[ 69] = 32'sh0692D04A;
        sine_table[ 70] = 32'sh06A9B20B; sine_table[ 71] = 32'sh06C0835B;
        sine_table[ 72] = 32'sh06D74402; sine_table[ 73] = 32'sh06EDF3C9;
        sine_table[ 74] = 32'sh07049276; sine_table[ 75] = 32'sh071B1FD2;
        sine_table[ 76] = 32'sh07319BA6; sine_table[ 77] = 32'sh074805BA;
        sine_table[ 78] = 32'sh075E5DD7; sine_table[ 79] = 32'sh0774A3C5;
        sine_table[ 80] = 32'sh078AD74E; sine_table[ 81] = 32'sh07A0F83B;
        sine_table[ 82] = 32'sh07B70655; sine_table[ 83] = 32'sh07CD0166;
        sine_table[ 84] = 32'sh07E2E937; sine_table[ 85] = 32'sh07F8BD93;
        sine_table[ 86] = 32'sh080E7E44; sine_table[ 87] = 32'sh08242B13;
        sine_table[ 88] = 32'sh0839C3CD; sine_table[ 89] = 32'sh084F483A;
        sine_table[ 90] = 32'sh0864B827; sine_table[ 91] = 32'sh087A135E;
        sine_table[ 92] = 32'sh088F59AA; sine_table[ 93] = 32'sh08A48AD8;
        sine_table[ 94] = 32'sh08B9A6B2; sine_table[ 95] = 32'sh08CEAD05;
        sine_table[ 96] = 32'sh08E39D9D; sine_table[ 97] = 32'sh08F87846;
        sine_table[ 98] = 32'sh090D3CCD; sine_table[ 99] = 32'sh0921EAFE;
        sine_table[100] = 32'sh093682A6; sine_table[101] = 32'sh094B0394;
        sine_table[102] = 32'sh095F6D93; sine_table[103] = 32'sh0973C072;
        sine_table[104] = 32'sh0987FBFE; sine_table[105] = 32'sh099C2007;
        sine_table[106] = 32'sh09B02C59; sine_table[107] = 32'sh09C420C3;
        sine_table[108] = 32'sh09D7FD15; sine_table[109] = 32'sh09EBC11C;
        sine_table[110] = 32'sh09FF6CAA; sine_table[111] = 32'sh0A12FF8C;
        sine_table[112] = 32'sh0A267993; sine_table[113] = 32'sh0A39DA8E;
        sine_table[114] = 32'sh0A4D224E; sine_table[115] = 32'sh0A6050A3;
        sine_table[116] = 32'sh0A73655E; sine_table[117] = 32'sh0A866050;
        sine_table[118] = 32'sh0A994149; sine_table[119] = 32'sh0AAC081C;
        sine_table[120] = 32'sh0ABEB49A; sine_table[121] = 32'sh0AD14695;
        sine_table[122] = 32'sh0AE3BDDF; sine_table[123] = 32'sh0AF61A4B;
        sine_table[124] = 32'sh0B085BAB; sine_table[125] = 32'sh0B1A81D2;
        sine_table[126] = 32'sh0B2C8C93; sine_table[127] = 32'sh0B3E7BC2;
        sine_table[128] = 32'sh0B504F33; sine_table[129] = 32'sh0B6206BA;
        sine_table[130] = 32'sh0B73A22A; sine_table[131] = 32'sh0B85215A;
        sine_table[132] = 32'sh0B96841C; sine_table[133] = 32'sh0BA7CA47;
        sine_table[134] = 32'sh0BB8F3B0; sine_table[135] = 32'sh0BCA002C;
        sine_table[136] = 32'sh0BDAEF91; sine_table[137] = 32'sh0BEBC1B6;
        sine_table[138] = 32'sh0BFC7672; sine_table[139] = 32'sh0C0D0D9A;
        sine_table[140] = 32'sh0C1D8706; sine_table[141] = 32'sh0C2DE28D;
        sine_table[142] = 32'sh0C3E2008; sine_table[143] = 32'sh0C4E3F4D;
        sine_table[144] = 32'sh0C5E4036; sine_table[145] = 32'sh0C6E229A;
        sine_table[146] = 32'sh0C7DE652; sine_table[147] = 32'sh0C8D8B38;
        sine_table[148] = 32'sh0C9D1125; sine_table[149] = 32'sh0CAC77F2;
        sine_table[150] = 32'sh0CBBBF7A; sine_table[151] = 32'sh0CCAE797;
        sine_table[152] = 32'sh0CD9F024; sine_table[153] = 32'sh0CE8D8FB;
        sine_table[154] = 32'sh0CF7A1F8; sine_table[155] = 32'sh0D064AF5;
        sine_table[156] = 32'sh0D14D3D0; sine_table[157] = 32'sh0D233C64;
        sine_table[158] = 32'sh0D31848E; sine_table[159] = 32'sh0D3FAC29;
        sine_table[160] = 32'sh0D4DB315; sine_table[161] = 32'sh0D5B992D;
        sine_table[162] = 32'sh0D695E4F; sine_table[163] = 32'sh0D77025A;
        sine_table[164] = 32'sh0D84852C; sine_table[165] = 32'sh0D91E6A4;
        sine_table[166] = 32'sh0D9F269F; sine_table[167] = 32'sh0DAC44FF;
        sine_table[168] = 32'sh0DB941A3; sine_table[169] = 32'sh0DC61C69;
        sine_table[170] = 32'sh0DD2D534; sine_table[171] = 32'sh0DDF6BE2;
        sine_table[172] = 32'sh0DEBE056; sine_table[173] = 32'sh0DF83271;
        sine_table[174] = 32'sh0E046213; sine_table[175] = 32'sh0E106F20;
        sine_table[176] = 32'sh0E1C5979; sine_table[177] = 32'sh0E282101;
        sine_table[178] = 32'sh0E33C59A; sine_table[179] = 32'sh0E3F4729;
        sine_table[180] = 32'sh0E4AA591; sine_table[181] = 32'sh0E55E0B5;
        sine_table[182] = 32'sh0E60F87A; sine_table[183] = 32'sh0E6BECC5;
        sine_table[184] = 32'sh0E76BD7A; sine_table[185] = 32'sh0E816A7F;
        sine_table[186] = 32'sh0E8BF3BA; sine_table[187] = 32'sh0E965910;
        sine_table[188] = 32'sh0EA09A69; sine_table[189] = 32'sh0EAAB7A9;
        sine_table[190] = 32'sh0EB4B0BA; sine_table[191] = 32'sh0EBE8581;
        sine_table[192] = 32'sh0EC835E8; sine_table[193] = 32'sh0ED1C1D5;
        sine_table[194] = 32'sh0EDB2931; sine_table[195] = 32'sh0EE46BE6;
        sine_table[196] = 32'sh0EED89DB; sine_table[197] = 32'sh0EF682FC;
        sine_table[198] = 32'sh0EFF5731; sine_table[199] = 32'sh0F080665;
        sine_table[200] = 32'sh0F109082; sine_table[201] = 32'sh0F18F574;
        sine_table[202] = 32'sh0F213526; sine_table[203] = 32'sh0F294F82;
        sine_table[204] = 32'sh0F314476; sine_table[205] = 32'sh0F3913EE;
        sine_table[206] = 32'sh0F40BDD6; sine_table[207] = 32'sh0F48421B;
        sine_table[208] = 32'sh0F4FA0AB; sine_table[209] = 32'sh0F56D974;
        sine_table[210] = 32'sh0F5DEC64; sine_table[211] = 32'sh0F64D96A;
        sine_table[212] = 32'sh0F6BA074; sine_table[213] = 32'sh0F724171;
        sine_table[214] = 32'sh0F78BC52; sine_table[215] = 32'sh0F7F1106;
        sine_table[216] = 32'sh0F853F7E; sine_table[217] = 32'sh0F8B47AA;
        sine_table[218] = 32'sh0F91297C; sine_table[219] = 32'sh0F96E4E5;
        sine_table[220] = 32'sh0F9C79D6; sine_table[221] = 32'sh0FA1E843;
        sine_table[222] = 32'sh0FA7301E; sine_table[223] = 32'sh0FAC5159;
        sine_table[224] = 32'sh0FB14BE8; sine_table[225] = 32'sh0FB61FBF;
        sine_table[226] = 32'sh0FBACCD2; sine_table[227] = 32'sh0FBF5315;
        sine_table[228] = 32'sh0FC3B27D; sine_table[229] = 32'sh0FC7EB00;
        sine_table[230] = 32'sh0FCBFC92; sine_table[231] = 32'sh0FCFE72B;
        sine_table[232] = 32'sh0FD3AAC0; sine_table[233] = 32'sh0FD74747;
        sine_table[234] = 32'sh0FDABCB9; sine_table[235] = 32'sh0FDE0B0C;
        sine_table[236] = 32'sh0FE13238; sine_table[237] = 32'sh0FE43236;
        sine_table[238] = 32'sh0FE70AFF; sine_table[239] = 32'sh0FE9BC8A;
        sine_table[240] = 32'sh0FEC46D2; sine_table[241] = 32'sh0FEEA9D0;
        sine_table[242] = 32'sh0FF0E57E; sine_table[243] = 32'sh0FF2F9D8;
        sine_table[244] = 32'sh0FF4E6D7; sine_table[245] = 32'sh0FF6AC76;
        sine_table[246] = 32'sh0FF84AB3; sine_table[247] = 32'sh0FF9C188;
        sine_table[248] = 32'sh0FFB10F2; sine_table[249] = 32'sh0FFC38ED;
        sine_table[250] = 32'sh0FFD3978; sine_table[251] = 32'sh0FFE128F;
        sine_table[252] = 32'sh0FFEC430; sine_table[253] = 32'sh0FFF4E5A;
        sine_table[254] = 32'sh0FFFB10B; sine_table[255] = 32'sh0FFFEC43;
    end

    // =========================================================
    // Stage 1: Reduce angle mod 2*pi, determine quadrant
    // =========================================================
    // We need angle in [0, 2*pi). For the quarter-wave approach:
    //   quadrant 0: [0, pi/2)      → table[idx]
    //   quadrant 1: [pi/2, pi)     → table[255-idx]
    //   quadrant 2: [pi, 3pi/2)    → -table[idx]
    //   quadrant 3: [3pi/2, 2pi)   → -table[255-idx]

    // Modular reduction: we use the fractional bits after dividing by 2*pi.
    // angle / (2*pi) gives us the fractional position in the cycle.
    // We approximate by using the upper bits of (angle * (1/(2*pi))).
    //
    // Simpler approach: since we only need 256 entries per quadrant,
    // we need 10 bits of phase (2 for quadrant + 8 for index).
    // phase = angle * 256*4 / (2*pi) = angle * 512/pi
    //
    // Even simpler: divide the angle space into 1024 steps.
    // phase[9:0] = (angle / (2*pi)) * 1024
    //
    // For Q4.28 with range [-8,+8), 2*pi ≈ 6.283
    // We compute: phase = (angle * PHASE_SCALE) >> 28
    // where PHASE_SCALE = 2^28 * 1024 / (2*pi) = 1024 / (2*pi) * 2^28
    //                   = 162.97... * 2^28 ≈ 43,741,844,462
    // That overflows 32 bits, so we use a different approach.
    //
    // Practical approach: extract phase from angle directly.
    // 2*pi in Q4.28 = 0x6487_ED51. We need (angle mod 2*pi) / (2*pi) * 1024.
    // Since we want to avoid division, we use bit manipulation:
    //
    // angle_pos = angle mod 2*pi (reduced to [0, 2*pi))
    // We know 2*pi ≈ 6.283, which fits in 3 integer bits of Q4.28.
    // A 10-bit phase index covering [0, 2*pi) means each step = 2*pi/1024.
    // 2*pi/1024 in Q4.28 = 0x6487_ED51 >> 10 = 0x19220 (approx)
    //
    // Alternative: multiply angle by reciprocal of 2*pi to get [0,1) fraction,
    // then take upper 10 bits as phase index.
    // 1/(2*pi) in Q4.28 = 0.15915... * 2^28 = 42,722,829 = 0x028B_E60D

    localparam signed [WIDTH-1:0] RECIP_TWO_PI = 32'sh028B_E60D;  // 1/(2*pi) in Q4.28

    reg [1:0]  quadrant_r;
    reg [7:0]  table_idx_r;
    reg        negate_r;
    reg        mirror_r;

    // Intermediate: multiply angle by 1/(2*pi) to get fractional turns
    // Result is Q4.28 representing fraction of full circle
    // We only need the fractional part (lower 28 bits) → 10 upper frac bits = phase
    wire signed [63:0] phase_product = angle * RECIP_TWO_PI;
    // phase_product is Q8.56. The fractional turn is in bits [55:0].
    // We want 10 bits of phase from the fractional part.
    // Bits [55:46] of product = upper 10 bits of fractional turn
    wire [9:0] phase_raw = phase_product[55:46];

    always @(posedge clk) begin
        quadrant_r <= phase_raw[9:8];
        // Mirror index in quadrants 1 and 3
        mirror_r   <= phase_raw[8];
        if (phase_raw[8])
            table_idx_r <= ~phase_raw[7:0];  // 255 - idx
        else
            table_idx_r <= phase_raw[7:0];
        // Negate in quadrants 2 and 3
        negate_r <= phase_raw[9];
    end

    // =========================================================
    // Stage 2: Table lookup and sign application
    // =========================================================
    wire signed [WIDTH-1:0] table_val = sine_table[table_idx_r];

    always @(posedge clk) begin
        if (negate_r)
            result <= -table_val;
        else
            result <= table_val;
    end

endmodule
