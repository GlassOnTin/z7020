initial begin
    weight_mem[0] = 32'h00000000;
    weight_mem[1] = 32'h00000000;
    weight_mem[2] = 32'h00000000;
    weight_mem[3] = 32'h00000000;
    weight_mem[4] = 32'h00000000;
    weight_mem[5] = 32'h00000000;
    weight_mem[6] = 32'h00000000;
    weight_mem[7] = 32'h00000000;
    weight_mem[8] = 32'h00000000;
    weight_mem[9] = 32'h00000000;
    weight_mem[10] = 32'h00000000;
    weight_mem[11] = 32'h00000000;
    weight_mem[12] = 32'h00000000;
    weight_mem[13] = 32'h00000000;
    weight_mem[14] = 32'h00000000;
    weight_mem[15] = 32'h00000000;
    weight_mem[16] = 32'h00000000;
    weight_mem[17] = 32'h00000000;
    weight_mem[18] = 32'h00000000;
    weight_mem[19] = 32'h00000000;
    weight_mem[20] = 32'h00000000;
    weight_mem[21] = 32'h00000000;
    weight_mem[22] = 32'h00000000;
    weight_mem[23] = 32'h00000000;
    weight_mem[24] = 32'h00000000;
    weight_mem[25] = 32'h00000000;
    weight_mem[26] = 32'h00000000;
    weight_mem[27] = 32'h00000000;
    weight_mem[28] = 32'h00000000;
    weight_mem[29] = 32'h00000000;
    weight_mem[30] = 32'h00000000;
    weight_mem[31] = 32'h00000000;
    weight_mem[32] = 32'h00000000;
    weight_mem[33] = 32'h00000000;
    weight_mem[34] = 32'h00000000;
    weight_mem[35] = 32'h00000000;
    weight_mem[36] = 32'h00000000;
    weight_mem[37] = 32'h00000000;
    weight_mem[38] = 32'h00000000;
    weight_mem[39] = 32'h00000000;
    weight_mem[40] = 32'h00000000;
    weight_mem[41] = 32'h00000000;
    weight_mem[42] = 32'h00000000;
    weight_mem[43] = 32'h00000000;
    weight_mem[44] = 32'h00000000;
    weight_mem[45] = 32'h00000000;
    weight_mem[46] = 32'h00000000;
    weight_mem[47] = 32'h00000000;
    weight_mem[48] = 32'h00000000;
    weight_mem[49] = 32'h00000000;
    weight_mem[50] = 32'h00000000;
    weight_mem[51] = 32'h00000000;
    weight_mem[52] = 32'h00000000;
    weight_mem[53] = 32'h00000000;
    weight_mem[54] = 32'h00000000;
    weight_mem[55] = 32'h00000000;
    weight_mem[56] = 32'h00000000;
    weight_mem[57] = 32'h00000000;
    weight_mem[58] = 32'h00000000;
    weight_mem[59] = 32'h00000000;
    weight_mem[60] = 32'h00000000;
    weight_mem[61] = 32'h00000000;
    weight_mem[62] = 32'h00000000;
    weight_mem[63] = 32'h00000000;
    weight_mem[64] = 32'h00000000;
    weight_mem[65] = 32'h00000000;
    weight_mem[66] = 32'h00000000;
    weight_mem[67] = 32'h00000000;
    weight_mem[68] = 32'h00000000;
    weight_mem[69] = 32'h00000000;
    weight_mem[70] = 32'h00000000;
    weight_mem[71] = 32'h00000000;
    weight_mem[72] = 32'h00000000;
    weight_mem[73] = 32'h00000000;
    weight_mem[74] = 32'h00000000;
    weight_mem[75] = 32'h00000000;
    weight_mem[76] = 32'h00000000;
    weight_mem[77] = 32'h00000000;
    weight_mem[78] = 32'h00000000;
    weight_mem[79] = 32'h00000000;
    weight_mem[80] = 32'h00000000;
    weight_mem[81] = 32'h00000000;
    weight_mem[82] = 32'h00000000;
    weight_mem[83] = 32'h00000000;
    weight_mem[84] = 32'h00000000;
    weight_mem[85] = 32'h00000000;
    weight_mem[86] = 32'h00000000;
    weight_mem[87] = 32'h00000000;
    weight_mem[88] = 32'h00000000;
    weight_mem[89] = 32'h00000000;
    weight_mem[90] = 32'h00000000;
    weight_mem[91] = 32'h00000000;
    weight_mem[92] = 32'h00000000;
    weight_mem[93] = 32'h00000000;
    weight_mem[94] = 32'h00000000;
    weight_mem[95] = 32'h00000000;
    weight_mem[96] = 32'h00000000;
    weight_mem[97] = 32'h00000000;
    weight_mem[98] = 32'h00000000;
    weight_mem[99] = 32'h00000000;
    weight_mem[100] = 32'h00000000;
    weight_mem[101] = 32'h00000000;
    weight_mem[102] = 32'h00000000;
    weight_mem[103] = 32'h00000000;
    weight_mem[104] = 32'h00000000;
    weight_mem[105] = 32'h00000000;
    weight_mem[106] = 32'h00000000;
    weight_mem[107] = 32'h00000000;
    weight_mem[108] = 32'h00000000;
    weight_mem[109] = 32'h00000000;
    weight_mem[110] = 32'h00000000;
    weight_mem[111] = 32'h00000000;
    weight_mem[112] = 32'h00000000;
    weight_mem[113] = 32'h00000000;
    weight_mem[114] = 32'h00000000;
    weight_mem[115] = 32'h00000000;
    weight_mem[116] = 32'h00000000;
    weight_mem[117] = 32'h00000000;
    weight_mem[118] = 32'h00000000;
    weight_mem[119] = 32'h00000000;
    weight_mem[120] = 32'h00000000;
    weight_mem[121] = 32'h00000000;
    weight_mem[122] = 32'h00000000;
    weight_mem[123] = 32'h00000000;
    weight_mem[124] = 32'h00000000;
    weight_mem[125] = 32'h00000000;
    weight_mem[126] = 32'h00000000;
    weight_mem[127] = 32'h00000000;
    weight_mem[128] = 32'h00000000;
    weight_mem[129] = 32'h00000000;
    weight_mem[130] = 32'h00000000;
    weight_mem[131] = 32'h00000000;
    weight_mem[132] = 32'h00000000;
    weight_mem[133] = 32'h00000000;
    weight_mem[134] = 32'h00000000;
    weight_mem[135] = 32'h00000000;
    weight_mem[136] = 32'h00000000;
    weight_mem[137] = 32'h00000000;
    weight_mem[138] = 32'h00000000;
    weight_mem[139] = 32'h00000000;
    weight_mem[140] = 32'h00000000;
    weight_mem[141] = 32'h00000000;
    weight_mem[142] = 32'h00000000;
    weight_mem[143] = 32'h00000000;
    weight_mem[144] = 32'h00000000;
    weight_mem[145] = 32'h00000000;
    weight_mem[146] = 32'h00000000;
    weight_mem[147] = 32'h00000000;
    weight_mem[148] = 32'h00000000;
    weight_mem[149] = 32'h00000000;
    weight_mem[150] = 32'h00000000;
    weight_mem[151] = 32'h00000000;
    weight_mem[152] = 32'h00000000;
    weight_mem[153] = 32'h00000000;
    weight_mem[154] = 32'h00000000;
    weight_mem[155] = 32'h00000000;
    weight_mem[156] = 32'h00000000;
    weight_mem[157] = 32'h00000000;
    weight_mem[158] = 32'h00000000;
    weight_mem[159] = 32'h00000000;
    weight_mem[160] = 32'h00000000;
    weight_mem[161] = 32'h00000000;
    weight_mem[162] = 32'h00000000;
    weight_mem[163] = 32'h00000000;
    weight_mem[164] = 32'h00000000;
    weight_mem[165] = 32'h00000000;
    weight_mem[166] = 32'h00000000;
    weight_mem[167] = 32'h00000000;
    weight_mem[168] = 32'h00000000;
    weight_mem[169] = 32'h00000000;
    weight_mem[170] = 32'h00000000;
    weight_mem[171] = 32'h00000000;
    weight_mem[172] = 32'h00000000;
    weight_mem[173] = 32'h00000000;
    weight_mem[174] = 32'h00000000;
    weight_mem[175] = 32'h00000000;
    weight_mem[176] = 32'h00000000;
    weight_mem[177] = 32'h00000000;
    weight_mem[178] = 32'h00000000;
    weight_mem[179] = 32'h00000000;
    weight_mem[180] = 32'h00000000;
    weight_mem[181] = 32'h00000000;
    weight_mem[182] = 32'h00000000;
    weight_mem[183] = 32'h00000000;
    weight_mem[184] = 32'h00000000;
    weight_mem[185] = 32'h00000000;
    weight_mem[186] = 32'h00000000;
    weight_mem[187] = 32'h00000000;
    weight_mem[188] = 32'h00000000;
    weight_mem[189] = 32'h00000000;
    weight_mem[190] = 32'h00000000;
    weight_mem[191] = 32'h00000000;
    weight_mem[192] = 32'h00000000;
    weight_mem[193] = 32'h00000000;
    weight_mem[194] = 32'h00000000;
    weight_mem[195] = 32'h00000000;
    weight_mem[196] = 32'h00000000;
    weight_mem[197] = 32'h00000000;
    weight_mem[198] = 32'h00000000;
    weight_mem[199] = 32'h00000000;
    weight_mem[200] = 32'h00000000;
    weight_mem[201] = 32'h00000000;
    weight_mem[202] = 32'h00000000;
    weight_mem[203] = 32'h00000000;
    weight_mem[204] = 32'h00000000;
    weight_mem[205] = 32'h00000000;
    weight_mem[206] = 32'h00000000;
    weight_mem[207] = 32'h00000000;
    weight_mem[208] = 32'h00000000;
    weight_mem[209] = 32'h00000000;
    weight_mem[210] = 32'h00000000;
    weight_mem[211] = 32'h00000000;
    weight_mem[212] = 32'h00000000;
    weight_mem[213] = 32'h00000000;
    weight_mem[214] = 32'h00000000;
    weight_mem[215] = 32'h00000000;
    weight_mem[216] = 32'h00000000;
    weight_mem[217] = 32'h00000000;
    weight_mem[218] = 32'h00000000;
    weight_mem[219] = 32'h00000000;
    weight_mem[220] = 32'h00000000;
    weight_mem[221] = 32'h00000000;
    weight_mem[222] = 32'h00000000;
    weight_mem[223] = 32'h00000000;
    weight_mem[224] = 32'h00000000;
    weight_mem[225] = 32'h00000000;
    weight_mem[226] = 32'h00000000;
    weight_mem[227] = 32'h00000000;
    weight_mem[228] = 32'h00000000;
    weight_mem[229] = 32'h00000000;
    weight_mem[230] = 32'h00000000;
    weight_mem[231] = 32'h00000000;
    weight_mem[232] = 32'h00000000;
    weight_mem[233] = 32'h00000000;
    weight_mem[234] = 32'h00000000;
    weight_mem[235] = 32'h00000000;
    weight_mem[236] = 32'h00000000;
    weight_mem[237] = 32'h00000000;
    weight_mem[238] = 32'h00000000;
    weight_mem[239] = 32'h00000000;
    weight_mem[240] = 32'h00000000;
    weight_mem[241] = 32'h00000000;
    weight_mem[242] = 32'h00000000;
    weight_mem[243] = 32'h00000000;
    weight_mem[244] = 32'h00000000;
    weight_mem[245] = 32'h00000000;
    weight_mem[246] = 32'h00000000;
    weight_mem[247] = 32'h00000000;
    weight_mem[248] = 32'h00000000;
    weight_mem[249] = 32'h00000000;
    weight_mem[250] = 32'h00000000;
    weight_mem[251] = 32'h00000000;
    weight_mem[252] = 32'h00000000;
    weight_mem[253] = 32'h00000000;
    weight_mem[254] = 32'h00000000;
    weight_mem[255] = 32'h00000000;
    weight_mem[256] = 32'h00000000;
    weight_mem[257] = 32'h00000000;
    weight_mem[258] = 32'h00000000;
    weight_mem[259] = 32'h00000000;
    weight_mem[260] = 32'h00000000;
    weight_mem[261] = 32'h00000000;
    weight_mem[262] = 32'h00000000;
    weight_mem[263] = 32'h00000000;
    weight_mem[264] = 32'h00000000;
    weight_mem[265] = 32'h00000000;
    weight_mem[266] = 32'h00000000;
    weight_mem[267] = 32'h00000000;
    weight_mem[268] = 32'h00000000;
    weight_mem[269] = 32'h00000000;
    weight_mem[270] = 32'h00000000;
    weight_mem[271] = 32'h00000000;
    weight_mem[272] = 32'h00000000;
    weight_mem[273] = 32'h00000000;
    weight_mem[274] = 32'h00000000;
    weight_mem[275] = 32'h00000000;
    weight_mem[276] = 32'h00000000;
    weight_mem[277] = 32'h00000000;
    weight_mem[278] = 32'h00000000;
    weight_mem[279] = 32'h00000000;
    weight_mem[280] = 32'h00000000;
    weight_mem[281] = 32'h00000000;
    weight_mem[282] = 32'h00000000;
    weight_mem[283] = 32'h00000000;
    weight_mem[284] = 32'h00000000;
    weight_mem[285] = 32'h00000000;
    weight_mem[286] = 32'h00000000;
    weight_mem[287] = 32'h00000000;
    weight_mem[288] = 32'h00000000;
    weight_mem[289] = 32'h00000000;
    weight_mem[290] = 32'h00000000;
    weight_mem[291] = 32'h00000000;
    weight_mem[292] = 32'h00000000;
    weight_mem[293] = 32'h00000000;
    weight_mem[294] = 32'h00000000;
    weight_mem[295] = 32'h00000000;
    weight_mem[296] = 32'h00000000;
    weight_mem[297] = 32'h00000000;
    weight_mem[298] = 32'h00000000;
    weight_mem[299] = 32'h00000000;
    weight_mem[300] = 32'h00000000;
    weight_mem[301] = 32'h00000000;
    weight_mem[302] = 32'h00000000;
    weight_mem[303] = 32'h00000000;
    weight_mem[304] = 32'h00000000;
    weight_mem[305] = 32'h00000000;
    weight_mem[306] = 32'h00000000;
    weight_mem[307] = 32'h00000000;
    weight_mem[308] = 32'h00000000;
    weight_mem[309] = 32'h00000000;
    weight_mem[310] = 32'h00000000;
    weight_mem[311] = 32'h00000000;
    weight_mem[312] = 32'h00000000;
    weight_mem[313] = 32'h00000000;
    weight_mem[314] = 32'h00000000;
    weight_mem[315] = 32'h00000000;
    weight_mem[316] = 32'h00000000;
    weight_mem[317] = 32'h00000000;
    weight_mem[318] = 32'h00000000;
    weight_mem[319] = 32'h00000000;
    weight_mem[320] = 32'h00000000;
    weight_mem[321] = 32'h00000000;
    weight_mem[322] = 32'h00000000;
    weight_mem[323] = 32'h00000000;
    weight_mem[324] = 32'h00000000;
    weight_mem[325] = 32'h00000000;
    weight_mem[326] = 32'h00000000;
    weight_mem[327] = 32'h00000000;
    weight_mem[328] = 32'h00000000;
    weight_mem[329] = 32'h00000000;
    weight_mem[330] = 32'h00000000;
    weight_mem[331] = 32'h00000000;
    weight_mem[332] = 32'h00000000;
    weight_mem[333] = 32'h00000000;
    weight_mem[334] = 32'h00000000;
    weight_mem[335] = 32'h00000000;
    weight_mem[336] = 32'h00000000;
    weight_mem[337] = 32'h00000000;
    weight_mem[338] = 32'h00000000;
    weight_mem[339] = 32'h00000000;
    weight_mem[340] = 32'h00000000;
    weight_mem[341] = 32'h00000000;
    weight_mem[342] = 32'h00000000;
    weight_mem[343] = 32'h00000000;
    weight_mem[344] = 32'h00000000;
    weight_mem[345] = 32'h00000000;
    weight_mem[346] = 32'h00000000;
    weight_mem[347] = 32'h00000000;
    weight_mem[348] = 32'h00000000;
    weight_mem[349] = 32'h00000000;
    weight_mem[350] = 32'h00000000;
    weight_mem[351] = 32'h00000000;
    weight_mem[352] = 32'h00000000;
    weight_mem[353] = 32'h00000000;
    weight_mem[354] = 32'h00000000;
    weight_mem[355] = 32'h00000000;
    weight_mem[356] = 32'h00000000;
    weight_mem[357] = 32'h00000000;
    weight_mem[358] = 32'h00000000;
    weight_mem[359] = 32'h00000000;
    weight_mem[360] = 32'h00000000;
    weight_mem[361] = 32'h00000000;
    weight_mem[362] = 32'h00000000;
    weight_mem[363] = 32'h00000000;
    weight_mem[364] = 32'h00000000;
    weight_mem[365] = 32'h00000000;
    weight_mem[366] = 32'h00000000;
    weight_mem[367] = 32'h00000000;
    weight_mem[368] = 32'h00000000;
    weight_mem[369] = 32'h00000000;
    weight_mem[370] = 32'h00000000;
    weight_mem[371] = 32'h00000000;
    weight_mem[372] = 32'h00000000;
    weight_mem[373] = 32'h00000000;
    weight_mem[374] = 32'h00000000;
    weight_mem[375] = 32'h00000000;
    weight_mem[376] = 32'h00000000;
    weight_mem[377] = 32'h00000000;
    weight_mem[378] = 32'h00000000;
    weight_mem[379] = 32'h00000000;
    weight_mem[380] = 32'h00000000;
    weight_mem[381] = 32'h00000000;
    weight_mem[382] = 32'h00000000;
    weight_mem[383] = 32'h00000000;
    weight_mem[384] = 32'h00000000;
    weight_mem[385] = 32'h00000000;
    weight_mem[386] = 32'h00000000;
    weight_mem[387] = 32'h00000000;
    weight_mem[388] = 32'h00000000;
    weight_mem[389] = 32'h00000000;
    weight_mem[390] = 32'h00000000;
    weight_mem[391] = 32'h00000000;
    weight_mem[392] = 32'h00000000;
    weight_mem[393] = 32'h00000000;
    weight_mem[394] = 32'h00000000;
    weight_mem[395] = 32'h00000000;
    weight_mem[396] = 32'h00000000;
    weight_mem[397] = 32'h00000000;
    weight_mem[398] = 32'h00000000;
    weight_mem[399] = 32'h00000000;
    weight_mem[400] = 32'h00000000;
    weight_mem[401] = 32'h00000000;
    weight_mem[402] = 32'h00000000;
    weight_mem[403] = 32'h00000000;
    weight_mem[404] = 32'h00000000;
    weight_mem[405] = 32'h00000000;
    weight_mem[406] = 32'h00000000;
    weight_mem[407] = 32'h00000000;
    weight_mem[408] = 32'h00000000;
    weight_mem[409] = 32'h00000000;
    weight_mem[410] = 32'h00000000;
    weight_mem[411] = 32'h00000000;
    weight_mem[412] = 32'h00000000;
    weight_mem[413] = 32'h00000000;
    weight_mem[414] = 32'h00000000;
    weight_mem[415] = 32'h00000000;
    weight_mem[416] = 32'h00000000;
    weight_mem[417] = 32'h00000000;
    weight_mem[418] = 32'h00000000;
    weight_mem[419] = 32'h00000000;
    weight_mem[420] = 32'h00000000;
    weight_mem[421] = 32'h00000000;
    weight_mem[422] = 32'h00000000;
    weight_mem[423] = 32'h00000000;
    weight_mem[424] = 32'h00000000;
    weight_mem[425] = 32'h00000000;
    weight_mem[426] = 32'h00000000;
    weight_mem[427] = 32'h00000000;
    weight_mem[428] = 32'h00000000;
    weight_mem[429] = 32'h00000000;
    weight_mem[430] = 32'h00000000;
    weight_mem[431] = 32'h00000000;
    weight_mem[432] = 32'h00000000;
    weight_mem[433] = 32'h00000000;
    weight_mem[434] = 32'h00000000;
    weight_mem[435] = 32'h00000000;
    weight_mem[436] = 32'h00000000;
    weight_mem[437] = 32'h00000000;
    weight_mem[438] = 32'h00000000;
    weight_mem[439] = 32'h00000000;
    weight_mem[440] = 32'h00000000;
    weight_mem[441] = 32'h00000000;
    weight_mem[442] = 32'h00000000;
    weight_mem[443] = 32'h00000000;
    weight_mem[444] = 32'h00000000;
    weight_mem[445] = 32'h00000000;
    weight_mem[446] = 32'h00000000;
    weight_mem[447] = 32'h00000000;
    weight_mem[448] = 32'h00000000;
    weight_mem[449] = 32'h00000000;
    weight_mem[450] = 32'h00000000;
    weight_mem[451] = 32'h00000000;
    weight_mem[452] = 32'h00000000;
    weight_mem[453] = 32'h00000000;
    weight_mem[454] = 32'h00000000;
    weight_mem[455] = 32'h00000000;
    weight_mem[456] = 32'h00000000;
    weight_mem[457] = 32'h00000000;
    weight_mem[458] = 32'h00000000;
    weight_mem[459] = 32'h00000000;
    weight_mem[460] = 32'h00000000;
    weight_mem[461] = 32'h00000000;
    weight_mem[462] = 32'h00000000;
    weight_mem[463] = 32'h00000000;
    weight_mem[464] = 32'h00000000;
    weight_mem[465] = 32'h00000000;
    weight_mem[466] = 32'h00000000;
    weight_mem[467] = 32'h00000000;
    weight_mem[468] = 32'h00000000;
    weight_mem[469] = 32'h00000000;
    weight_mem[470] = 32'h00000000;
    weight_mem[471] = 32'h00000000;
    weight_mem[472] = 32'h00000000;
    weight_mem[473] = 32'h00000000;
    weight_mem[474] = 32'h00000000;
    weight_mem[475] = 32'h00000000;
    weight_mem[476] = 32'h00000000;
    weight_mem[477] = 32'h00000000;
    weight_mem[478] = 32'h00000000;
    weight_mem[479] = 32'h00000000;
    weight_mem[480] = 32'h00000000;
    weight_mem[481] = 32'h00000000;
    weight_mem[482] = 32'h00000000;
    weight_mem[483] = 32'h00000000;
    weight_mem[484] = 32'h00000000;
    weight_mem[485] = 32'h00000000;
    weight_mem[486] = 32'h00000000;
    weight_mem[487] = 32'h00000000;
    weight_mem[488] = 32'h00000000;
    weight_mem[489] = 32'h00000000;
    weight_mem[490] = 32'h00000000;
    weight_mem[491] = 32'h00000000;
    weight_mem[492] = 32'h00000000;
    weight_mem[493] = 32'h00000000;
    weight_mem[494] = 32'h00000000;
    weight_mem[495] = 32'h00000000;
    weight_mem[496] = 32'h00000000;
    weight_mem[497] = 32'h00000000;
    weight_mem[498] = 32'h00000000;
    weight_mem[499] = 32'h00000000;
    weight_mem[500] = 32'h00000000;
    weight_mem[501] = 32'h00000000;
    weight_mem[502] = 32'h00000000;
    weight_mem[503] = 32'h00000000;
    weight_mem[504] = 32'h00000000;
    weight_mem[505] = 32'h00000000;
    weight_mem[506] = 32'h00000000;
    weight_mem[507] = 32'h00000000;
    weight_mem[508] = 32'h00000000;
    weight_mem[509] = 32'h00000000;
    weight_mem[510] = 32'h00000000;
    weight_mem[511] = 32'h00000000;
    weight_mem[512] = 32'h00000000;
    weight_mem[513] = 32'h00000000;
    weight_mem[514] = 32'h00000000;
    weight_mem[515] = 32'h00000000;
    weight_mem[516] = 32'h00000000;
    weight_mem[517] = 32'h00000000;
    weight_mem[518] = 32'h00000000;
    weight_mem[519] = 32'h00000000;
    weight_mem[520] = 32'h00000000;
    weight_mem[521] = 32'h00000000;
    weight_mem[522] = 32'h00000000;
    weight_mem[523] = 32'h00000000;
    weight_mem[524] = 32'h00000000;
    weight_mem[525] = 32'h00000000;
    weight_mem[526] = 32'h00000000;
    weight_mem[527] = 32'h00000000;
    weight_mem[528] = 32'h00000000;
    weight_mem[529] = 32'h00000000;
    weight_mem[530] = 32'h00000000;
    weight_mem[531] = 32'h00000000;
    weight_mem[532] = 32'h00000000;
    weight_mem[533] = 32'h00000000;
    weight_mem[534] = 32'h00000000;
    weight_mem[535] = 32'h00000000;
    weight_mem[536] = 32'h00000000;
    weight_mem[537] = 32'h00000000;
    weight_mem[538] = 32'h00000000;
    weight_mem[539] = 32'h00000000;
    weight_mem[540] = 32'h00000000;
    weight_mem[541] = 32'h00000000;
    weight_mem[542] = 32'h00000000;
    weight_mem[543] = 32'h00000000;
    weight_mem[544] = 32'h00000000;
    weight_mem[545] = 32'h00000000;
    weight_mem[546] = 32'h00000000;
    weight_mem[547] = 32'h00000000;
    weight_mem[548] = 32'h00000000;
    weight_mem[549] = 32'h00000000;
    weight_mem[550] = 32'h00000000;
    weight_mem[551] = 32'h00000000;
    weight_mem[552] = 32'h00000000;
    weight_mem[553] = 32'h00000000;
    weight_mem[554] = 32'h00000000;
    weight_mem[555] = 32'h00000000;
    weight_mem[556] = 32'h00000000;
    weight_mem[557] = 32'h00000000;
    weight_mem[558] = 32'h00000000;
    weight_mem[559] = 32'h00000000;
    weight_mem[560] = 32'h00000000;
    weight_mem[561] = 32'h00000000;
    weight_mem[562] = 32'h00000000;
    weight_mem[563] = 32'h00000000;
    weight_mem[564] = 32'h00000000;
    weight_mem[565] = 32'h00000000;
    weight_mem[566] = 32'h00000000;
    weight_mem[567] = 32'h00000000;
    weight_mem[568] = 32'h00000000;
    weight_mem[569] = 32'h00000000;
    weight_mem[570] = 32'h00000000;
    weight_mem[571] = 32'h00000000;
    weight_mem[572] = 32'h00000000;
    weight_mem[573] = 32'h00000000;
    weight_mem[574] = 32'h00000000;
    weight_mem[575] = 32'h00000000;
    weight_mem[576] = 32'h00000000;
    weight_mem[577] = 32'h00000000;
    weight_mem[578] = 32'h00000000;
    weight_mem[579] = 32'h00000000;
    weight_mem[580] = 32'h00000000;
    weight_mem[581] = 32'h00000000;
    weight_mem[582] = 32'h00000000;
    weight_mem[583] = 32'h00000000;
    weight_mem[584] = 32'h00000000;
    weight_mem[585] = 32'h00000000;
    weight_mem[586] = 32'h00000000;
    weight_mem[587] = 32'h00000000;
    weight_mem[588] = 32'h00000000;
    weight_mem[589] = 32'h00000000;
    weight_mem[590] = 32'h00000000;
    weight_mem[591] = 32'h00000000;
    weight_mem[592] = 32'h00000000;
    weight_mem[593] = 32'h00000000;
    weight_mem[594] = 32'h00000000;
    weight_mem[595] = 32'h00000000;
    weight_mem[596] = 32'h00000000;
    weight_mem[597] = 32'h00000000;
    weight_mem[598] = 32'h00000000;
    weight_mem[599] = 32'h00000000;
    weight_mem[600] = 32'h00000000;
    weight_mem[601] = 32'h00000000;
    weight_mem[602] = 32'h00000000;
    weight_mem[603] = 32'h00000000;
    weight_mem[604] = 32'h00000000;
    weight_mem[605] = 32'h00000000;
    weight_mem[606] = 32'h00000000;
    weight_mem[607] = 32'h00000000;
    weight_mem[608] = 32'h00000000;
    weight_mem[609] = 32'h00000000;
    weight_mem[610] = 32'h00000000;
    weight_mem[611] = 32'h00000000;
    weight_mem[612] = 32'h00000000;
    weight_mem[613] = 32'h00000000;
    weight_mem[614] = 32'h00000000;
    weight_mem[615] = 32'h00000000;
    weight_mem[616] = 32'h00000000;
    weight_mem[617] = 32'h00000000;
    weight_mem[618] = 32'h00000000;
    weight_mem[619] = 32'h00000000;
    weight_mem[620] = 32'h00000000;
    weight_mem[621] = 32'h00000000;
    weight_mem[622] = 32'h00000000;
    weight_mem[623] = 32'h00000000;
    weight_mem[624] = 32'h00000000;
    weight_mem[625] = 32'h00000000;
    weight_mem[626] = 32'h00000000;
    weight_mem[627] = 32'h00000000;
    weight_mem[628] = 32'h00000000;
    weight_mem[629] = 32'h00000000;
    weight_mem[630] = 32'h00000000;
    weight_mem[631] = 32'h00000000;
    weight_mem[632] = 32'h00000000;
    weight_mem[633] = 32'h00000000;
    weight_mem[634] = 32'h00000000;
    weight_mem[635] = 32'h00000000;
    weight_mem[636] = 32'h00000000;
    weight_mem[637] = 32'h00000000;
    weight_mem[638] = 32'h00000000;
    weight_mem[639] = 32'h00000000;
    weight_mem[640] = 32'h00000000;
    weight_mem[641] = 32'h00000000;
    weight_mem[642] = 32'h00000000;
    weight_mem[643] = 32'h00000000;
    weight_mem[644] = 32'h00000000;
    weight_mem[645] = 32'h00000000;
    weight_mem[646] = 32'h00000000;
    weight_mem[647] = 32'h00000000;
    weight_mem[648] = 32'h00000000;
    weight_mem[649] = 32'h00000000;
    weight_mem[650] = 32'h00000000;
    weight_mem[651] = 32'h00000000;
    weight_mem[652] = 32'h00000000;
    weight_mem[653] = 32'h00000000;
    weight_mem[654] = 32'h00000000;
    weight_mem[655] = 32'h00000000;
    weight_mem[656] = 32'h00000000;
    weight_mem[657] = 32'h00000000;
    weight_mem[658] = 32'h00000000;
    weight_mem[659] = 32'h00000000;
    weight_mem[660] = 32'h00000000;
    weight_mem[661] = 32'h00000000;
    weight_mem[662] = 32'h00000000;
    weight_mem[663] = 32'h00000000;
    weight_mem[664] = 32'h00000000;
    weight_mem[665] = 32'h00000000;
    weight_mem[666] = 32'h00000000;
    weight_mem[667] = 32'h00000000;
    weight_mem[668] = 32'h00000000;
    weight_mem[669] = 32'h00000000;
    weight_mem[670] = 32'h00000000;
    weight_mem[671] = 32'h00000000;
    weight_mem[672] = 32'h00000000;
    weight_mem[673] = 32'h00000000;
    weight_mem[674] = 32'h00000000;
    weight_mem[675] = 32'h00000000;
    weight_mem[676] = 32'h00000000;
    weight_mem[677] = 32'h00000000;
    weight_mem[678] = 32'h00000000;
    weight_mem[679] = 32'h00000000;
    weight_mem[680] = 32'h00000000;
    weight_mem[681] = 32'h00000000;
    weight_mem[682] = 32'h00000000;
    weight_mem[683] = 32'h00000000;
    weight_mem[684] = 32'h00000000;
    weight_mem[685] = 32'h00000000;
    weight_mem[686] = 32'h00000000;
    weight_mem[687] = 32'h00000000;
    weight_mem[688] = 32'h00000000;
    weight_mem[689] = 32'h00000000;
    weight_mem[690] = 32'h00000000;
    weight_mem[691] = 32'h00000000;
    weight_mem[692] = 32'h00000000;
    weight_mem[693] = 32'h00000000;
    weight_mem[694] = 32'h00000000;
    weight_mem[695] = 32'h00000000;
    weight_mem[696] = 32'h00000000;
    weight_mem[697] = 32'h00000000;
    weight_mem[698] = 32'h00000000;
    weight_mem[699] = 32'h00000000;
    weight_mem[700] = 32'h00000000;
    weight_mem[701] = 32'h00000000;
    weight_mem[702] = 32'h00000000;
    weight_mem[703] = 32'h00000000;
    weight_mem[704] = 32'h00000000;
    weight_mem[705] = 32'h00000000;
    weight_mem[706] = 32'h00000000;
    weight_mem[707] = 32'h00000000;
    weight_mem[708] = 32'h00000000;
    weight_mem[709] = 32'h00000000;
    weight_mem[710] = 32'h00000000;
    weight_mem[711] = 32'h00000000;
    weight_mem[712] = 32'h00000000;
    weight_mem[713] = 32'h00000000;
    weight_mem[714] = 32'h00000000;
    weight_mem[715] = 32'h00000000;
    weight_mem[716] = 32'h00000000;
    weight_mem[717] = 32'h00000000;
    weight_mem[718] = 32'h00000000;
    weight_mem[719] = 32'h00000000;
    weight_mem[720] = 32'h00000000;
    weight_mem[721] = 32'h00000000;
    weight_mem[722] = 32'h00000000;
    weight_mem[723] = 32'h00000000;
    weight_mem[724] = 32'h00000000;
    weight_mem[725] = 32'h00000000;
    weight_mem[726] = 32'h00000000;
    weight_mem[727] = 32'h00000000;
    weight_mem[728] = 32'h00000000;
    weight_mem[729] = 32'h00000000;
    weight_mem[730] = 32'h00000000;
    weight_mem[731] = 32'h00000000;
    weight_mem[732] = 32'h00000000;
    weight_mem[733] = 32'h00000000;
    weight_mem[734] = 32'h00000000;
    weight_mem[735] = 32'h00000000;
    weight_mem[736] = 32'h00000000;
    weight_mem[737] = 32'h00000000;
    weight_mem[738] = 32'h00000000;
    weight_mem[739] = 32'h00000000;
    weight_mem[740] = 32'h00000000;
    weight_mem[741] = 32'h00000000;
    weight_mem[742] = 32'h00000000;
    weight_mem[743] = 32'h00000000;
    weight_mem[744] = 32'h00000000;
    weight_mem[745] = 32'h00000000;
    weight_mem[746] = 32'h00000000;
    weight_mem[747] = 32'h00000000;
    weight_mem[748] = 32'h00000000;
    weight_mem[749] = 32'h00000000;
    weight_mem[750] = 32'h00000000;
    weight_mem[751] = 32'h00000000;
    weight_mem[752] = 32'h00000000;
    weight_mem[753] = 32'h00000000;
    weight_mem[754] = 32'h00000000;
    weight_mem[755] = 32'h00000000;
    weight_mem[756] = 32'h00000000;
    weight_mem[757] = 32'h00000000;
    weight_mem[758] = 32'h00000000;
    weight_mem[759] = 32'h00000000;
    weight_mem[760] = 32'h00000000;
    weight_mem[761] = 32'h00000000;
    weight_mem[762] = 32'h00000000;
    weight_mem[763] = 32'h00000000;
    weight_mem[764] = 32'h00000000;
    weight_mem[765] = 32'h00000000;
    weight_mem[766] = 32'h00000000;
    weight_mem[767] = 32'h00000000;
    weight_mem[768] = 32'h00000000;
    weight_mem[769] = 32'h00000000;
    weight_mem[770] = 32'h00000000;
    weight_mem[771] = 32'h00000000;
    weight_mem[772] = 32'h00000000;
    weight_mem[773] = 32'h00000000;
    weight_mem[774] = 32'h00000000;
    weight_mem[775] = 32'h00000000;
    weight_mem[776] = 32'h00000000;
    weight_mem[777] = 32'h00000000;
    weight_mem[778] = 32'h00000000;
    weight_mem[779] = 32'h00000000;
    weight_mem[780] = 32'h00000000;
    weight_mem[781] = 32'h00000000;
    weight_mem[782] = 32'h00000000;
    weight_mem[783] = 32'h00000000;
    weight_mem[784] = 32'h00000000;
    weight_mem[785] = 32'h00000000;
    weight_mem[786] = 32'h00000000;
    weight_mem[787] = 32'h00000000;
    weight_mem[788] = 32'h00000000;
    weight_mem[789] = 32'h00000000;
    weight_mem[790] = 32'h00000000;
    weight_mem[791] = 32'h00000000;
    weight_mem[792] = 32'h00000000;
    weight_mem[793] = 32'h00000000;
    weight_mem[794] = 32'h00000000;
    weight_mem[795] = 32'h00000000;
    weight_mem[796] = 32'h00000000;
    weight_mem[797] = 32'h00000000;
    weight_mem[798] = 32'h00000000;
    weight_mem[799] = 32'h00000000;
    weight_mem[800] = 32'h00000000;
    weight_mem[801] = 32'h00000000;
    weight_mem[802] = 32'h00000000;
    weight_mem[803] = 32'h00000000;
    weight_mem[804] = 32'h00000000;
    weight_mem[805] = 32'h00000000;
    weight_mem[806] = 32'h00000000;
    weight_mem[807] = 32'h00000000;
    weight_mem[808] = 32'h00000000;
    weight_mem[809] = 32'h00000000;
    weight_mem[810] = 32'h00000000;
    weight_mem[811] = 32'h00000000;
    weight_mem[812] = 32'h00000000;
    weight_mem[813] = 32'h00000000;
    weight_mem[814] = 32'h00000000;
    weight_mem[815] = 32'h00000000;
    weight_mem[816] = 32'h00000000;
    weight_mem[817] = 32'h00000000;
    weight_mem[818] = 32'h00000000;
    weight_mem[819] = 32'h00000000;
    weight_mem[820] = 32'h00000000;
    weight_mem[821] = 32'h00000000;
    weight_mem[822] = 32'h00000000;
    weight_mem[823] = 32'h00000000;
    weight_mem[824] = 32'h00000000;
    weight_mem[825] = 32'h00000000;
    weight_mem[826] = 32'h00000000;
    weight_mem[827] = 32'h00000000;
    weight_mem[828] = 32'h00000000;
    weight_mem[829] = 32'h00000000;
    weight_mem[830] = 32'h00000000;
    weight_mem[831] = 32'h00000000;
    weight_mem[832] = 32'h00000000;
    weight_mem[833] = 32'h00000000;
    weight_mem[834] = 32'h00000000;
    weight_mem[835] = 32'h00000000;
    weight_mem[836] = 32'h00000000;
    weight_mem[837] = 32'h00000000;
    weight_mem[838] = 32'h00000000;
    weight_mem[839] = 32'h00000000;
    weight_mem[840] = 32'h00000000;
    weight_mem[841] = 32'h00000000;
    weight_mem[842] = 32'h00000000;
    weight_mem[843] = 32'h00000000;
    weight_mem[844] = 32'h00000000;
    weight_mem[845] = 32'h00000000;
    weight_mem[846] = 32'h00000000;
    weight_mem[847] = 32'h00000000;
    weight_mem[848] = 32'h00000000;
    weight_mem[849] = 32'h00000000;
    weight_mem[850] = 32'h00000000;
    weight_mem[851] = 32'h00000000;
    weight_mem[852] = 32'h00000000;
    weight_mem[853] = 32'h00000000;
    weight_mem[854] = 32'h00000000;
    weight_mem[855] = 32'h00000000;
    weight_mem[856] = 32'h00000000;
    weight_mem[857] = 32'h00000000;
    weight_mem[858] = 32'h00000000;
    weight_mem[859] = 32'h00000000;
    weight_mem[860] = 32'h00000000;
    weight_mem[861] = 32'h00000000;
    weight_mem[862] = 32'h00000000;
    weight_mem[863] = 32'h00000000;
    weight_mem[864] = 32'h00000000;
    weight_mem[865] = 32'h00000000;
    weight_mem[866] = 32'h00000000;
    weight_mem[867] = 32'h00000000;
    weight_mem[868] = 32'h00000000;
    weight_mem[869] = 32'h00000000;
    weight_mem[870] = 32'h00000000;
    weight_mem[871] = 32'h00000000;
    weight_mem[872] = 32'h00000000;
    weight_mem[873] = 32'h00000000;
    weight_mem[874] = 32'h00000000;
    weight_mem[875] = 32'h00000000;
    weight_mem[876] = 32'h00000000;
    weight_mem[877] = 32'h00000000;
    weight_mem[878] = 32'h00000000;
    weight_mem[879] = 32'h00000000;
    weight_mem[880] = 32'h00000000;
    weight_mem[881] = 32'h00000000;
    weight_mem[882] = 32'h00000000;
    weight_mem[883] = 32'h00000000;
    weight_mem[884] = 32'h00000000;
    weight_mem[885] = 32'h00000000;
    weight_mem[886] = 32'h00000000;
    weight_mem[887] = 32'h00000000;
    weight_mem[888] = 32'h00000000;
    weight_mem[889] = 32'h00000000;
    weight_mem[890] = 32'h00000000;
    weight_mem[891] = 32'h00000000;
    weight_mem[892] = 32'h00000000;
    weight_mem[893] = 32'h00000000;
    weight_mem[894] = 32'h00000000;
    weight_mem[895] = 32'h00000000;
    weight_mem[896] = 32'h00000000;
    weight_mem[897] = 32'h00000000;
    weight_mem[898] = 32'h00000000;
    weight_mem[899] = 32'h00000000;
    weight_mem[900] = 32'h00000000;
    weight_mem[901] = 32'h00000000;
    weight_mem[902] = 32'h00000000;
    weight_mem[903] = 32'h00000000;
    weight_mem[904] = 32'h00000000;
    weight_mem[905] = 32'h00000000;
    weight_mem[906] = 32'h00000000;
    weight_mem[907] = 32'h00000000;
    weight_mem[908] = 32'h00000000;
    weight_mem[909] = 32'h00000000;
    weight_mem[910] = 32'h00000000;
    weight_mem[911] = 32'h00000000;
    weight_mem[912] = 32'h00000000;
    weight_mem[913] = 32'h00000000;
    weight_mem[914] = 32'h00000000;
    weight_mem[915] = 32'h00000000;
    weight_mem[916] = 32'h00000000;
    weight_mem[917] = 32'h00000000;
    weight_mem[918] = 32'h00000000;
    weight_mem[919] = 32'h00000000;
    weight_mem[920] = 32'h00000000;
    weight_mem[921] = 32'h00000000;
    weight_mem[922] = 32'h00000000;
    weight_mem[923] = 32'h00000000;
    weight_mem[924] = 32'h00000000;
    weight_mem[925] = 32'h00000000;
    weight_mem[926] = 32'h00000000;
    weight_mem[927] = 32'h00000000;
    weight_mem[928] = 32'h00000000;
    weight_mem[929] = 32'h00000000;
    weight_mem[930] = 32'h00000000;
    weight_mem[931] = 32'h00000000;
    weight_mem[932] = 32'h00000000;
    weight_mem[933] = 32'h00000000;
    weight_mem[934] = 32'h00000000;
    weight_mem[935] = 32'h00000000;
    weight_mem[936] = 32'h00000000;
    weight_mem[937] = 32'h00000000;
    weight_mem[938] = 32'h00000000;
    weight_mem[939] = 32'h00000000;
    weight_mem[940] = 32'h00000000;
    weight_mem[941] = 32'h00000000;
    weight_mem[942] = 32'h00000000;
    weight_mem[943] = 32'h00000000;
    weight_mem[944] = 32'h00000000;
    weight_mem[945] = 32'h00000000;
    weight_mem[946] = 32'h00000000;
    weight_mem[947] = 32'h00000000;
    weight_mem[948] = 32'h00000000;
    weight_mem[949] = 32'h00000000;
    weight_mem[950] = 32'h00000000;
    weight_mem[951] = 32'h00000000;
    weight_mem[952] = 32'h00000000;
    weight_mem[953] = 32'h00000000;
    weight_mem[954] = 32'h00000000;
    weight_mem[955] = 32'h00000000;
    weight_mem[956] = 32'h00000000;
    weight_mem[957] = 32'h00000000;
    weight_mem[958] = 32'h00000000;
    weight_mem[959] = 32'h00000000;
    weight_mem[960] = 32'h00000000;
    weight_mem[961] = 32'h00000000;
    weight_mem[962] = 32'h00000000;
    weight_mem[963] = 32'h00000000;
    weight_mem[964] = 32'h00000000;
    weight_mem[965] = 32'h00000000;
    weight_mem[966] = 32'h00000000;
    weight_mem[967] = 32'h00000000;
    weight_mem[968] = 32'h00000000;
    weight_mem[969] = 32'h00000000;
    weight_mem[970] = 32'h00000000;
    weight_mem[971] = 32'h00000000;
    weight_mem[972] = 32'h00000000;
    weight_mem[973] = 32'h00000000;
    weight_mem[974] = 32'h00000000;
    weight_mem[975] = 32'h00000000;
    weight_mem[976] = 32'h00000000;
    weight_mem[977] = 32'h00000000;
    weight_mem[978] = 32'h00000000;
    weight_mem[979] = 32'h00000000;
    weight_mem[980] = 32'h00000000;
    weight_mem[981] = 32'h00000000;
    weight_mem[982] = 32'h00000000;
    weight_mem[983] = 32'h00000000;
    weight_mem[984] = 32'h00000000;
    weight_mem[985] = 32'h00000000;
    weight_mem[986] = 32'h00000000;
    weight_mem[987] = 32'h00000000;
    weight_mem[988] = 32'h00000000;
    weight_mem[989] = 32'h00000000;
    weight_mem[990] = 32'h00000000;
    weight_mem[991] = 32'h00000000;
    weight_mem[992] = 32'h00000000;
    weight_mem[993] = 32'h00000000;
    weight_mem[994] = 32'h00000000;
    weight_mem[995] = 32'h00000000;
    weight_mem[996] = 32'h00000000;
    weight_mem[997] = 32'h00000000;
    weight_mem[998] = 32'h00000000;
    weight_mem[999] = 32'h00000000;
    weight_mem[1000] = 32'h00000000;
    weight_mem[1001] = 32'h00000000;
    weight_mem[1002] = 32'h00000000;
    weight_mem[1003] = 32'h00000000;
    weight_mem[1004] = 32'h00000000;
    weight_mem[1005] = 32'h00000000;
    weight_mem[1006] = 32'h00000000;
    weight_mem[1007] = 32'h00000000;
    weight_mem[1008] = 32'h00000000;
    weight_mem[1009] = 32'h00000000;
    weight_mem[1010] = 32'h00000000;
    weight_mem[1011] = 32'h00000000;
    weight_mem[1012] = 32'h00000000;
    weight_mem[1013] = 32'h00000000;
    weight_mem[1014] = 32'h00000000;
    weight_mem[1015] = 32'h00000000;
    weight_mem[1016] = 32'h00000000;
    weight_mem[1017] = 32'h00000000;
    weight_mem[1018] = 32'h00000000;
    weight_mem[1019] = 32'h00000000;
    weight_mem[1020] = 32'h00000000;
    weight_mem[1021] = 32'h00000000;
    weight_mem[1022] = 32'h00000000;
    weight_mem[1023] = 32'h00000000;
    weight_mem[1024] = 32'h00000000;
    weight_mem[1025] = 32'h00000000;
    weight_mem[1026] = 32'h00000000;
    weight_mem[1027] = 32'h00000000;
    weight_mem[1028] = 32'h00000000;
    weight_mem[1029] = 32'h00000000;
    weight_mem[1030] = 32'h00000000;
    weight_mem[1031] = 32'h00000000;
    weight_mem[1032] = 32'h00000000;
    weight_mem[1033] = 32'h00000000;
    weight_mem[1034] = 32'h00000000;
    weight_mem[1035] = 32'h00000000;
    weight_mem[1036] = 32'h00000000;
    weight_mem[1037] = 32'h00000000;
    weight_mem[1038] = 32'h00000000;
    weight_mem[1039] = 32'h00000000;
    weight_mem[1040] = 32'h00000000;
    weight_mem[1041] = 32'h00000000;
    weight_mem[1042] = 32'h00000000;
    weight_mem[1043] = 32'h00000000;
    weight_mem[1044] = 32'h00000000;
    weight_mem[1045] = 32'h00000000;
    weight_mem[1046] = 32'h00000000;
    weight_mem[1047] = 32'h00000000;
    weight_mem[1048] = 32'h00000000;
    weight_mem[1049] = 32'h00000000;
    weight_mem[1050] = 32'h00000000;
    weight_mem[1051] = 32'h00000000;
    weight_mem[1052] = 32'h00000000;
    weight_mem[1053] = 32'h00000000;
    weight_mem[1054] = 32'h00000000;
    weight_mem[1055] = 32'h00000000;
    weight_mem[1056] = 32'h00000000;
    weight_mem[1057] = 32'h00000000;
    weight_mem[1058] = 32'h00000000;
    weight_mem[1059] = 32'h00000000;
    weight_mem[1060] = 32'h00000000;
    weight_mem[1061] = 32'h00000000;
    weight_mem[1062] = 32'h00000000;
    weight_mem[1063] = 32'h00000000;
    weight_mem[1064] = 32'h00000000;
    weight_mem[1065] = 32'h00000000;
    weight_mem[1066] = 32'h00000000;
    weight_mem[1067] = 32'h00000000;
    weight_mem[1068] = 32'h00000000;
    weight_mem[1069] = 32'h00000000;
    weight_mem[1070] = 32'h00000000;
    weight_mem[1071] = 32'h00000000;
    weight_mem[1072] = 32'h00000000;
    weight_mem[1073] = 32'h00000000;
    weight_mem[1074] = 32'h00000000;
    weight_mem[1075] = 32'h00000000;
    weight_mem[1076] = 32'h00000000;
    weight_mem[1077] = 32'h00000000;
    weight_mem[1078] = 32'h00000000;
    weight_mem[1079] = 32'h00000000;
    weight_mem[1080] = 32'h00000000;
    weight_mem[1081] = 32'h00000000;
    weight_mem[1082] = 32'h00000000;
    weight_mem[1083] = 32'h00000000;
    weight_mem[1084] = 32'h00000000;
    weight_mem[1085] = 32'h00000000;
    weight_mem[1086] = 32'h00000000;
    weight_mem[1087] = 32'h00000000;
    weight_mem[1088] = 32'h00000000;
    weight_mem[1089] = 32'h00000000;
    weight_mem[1090] = 32'h00000000;
    weight_mem[1091] = 32'h00000000;
    weight_mem[1092] = 32'h00000000;
    weight_mem[1093] = 32'h00000000;
    weight_mem[1094] = 32'h00000000;
    weight_mem[1095] = 32'h00000000;
    weight_mem[1096] = 32'h00000000;
    weight_mem[1097] = 32'h00000000;
    weight_mem[1098] = 32'h00000000;
    weight_mem[1099] = 32'h00000000;
    weight_mem[1100] = 32'h00000000;
    weight_mem[1101] = 32'h00000000;
    weight_mem[1102] = 32'h00000000;
    weight_mem[1103] = 32'h00000000;
    weight_mem[1104] = 32'h00000000;
    weight_mem[1105] = 32'h00000000;
    weight_mem[1106] = 32'h00000000;
    weight_mem[1107] = 32'h00000000;
    weight_mem[1108] = 32'h00000000;
    weight_mem[1109] = 32'h00000000;
    weight_mem[1110] = 32'h00000000;
    weight_mem[1111] = 32'h00000000;
    weight_mem[1112] = 32'h00000000;
    weight_mem[1113] = 32'h00000000;
    weight_mem[1114] = 32'h00000000;
    weight_mem[1115] = 32'h00000000;
    weight_mem[1116] = 32'h00000000;
    weight_mem[1117] = 32'h00000000;
    weight_mem[1118] = 32'h00000000;
    weight_mem[1119] = 32'h00000000;
    weight_mem[1120] = 32'h00000000;
    weight_mem[1121] = 32'h00000000;
    weight_mem[1122] = 32'h00000000;
    weight_mem[1123] = 32'h00000000;
    weight_mem[1124] = 32'h00000000;
    weight_mem[1125] = 32'h00000000;
    weight_mem[1126] = 32'h00000000;
    weight_mem[1127] = 32'h00000000;
    weight_mem[1128] = 32'h00000000;
    weight_mem[1129] = 32'h00000000;
    weight_mem[1130] = 32'h00000000;
    weight_mem[1131] = 32'h00000000;
    weight_mem[1132] = 32'h00000000;
    weight_mem[1133] = 32'h00000000;
    weight_mem[1134] = 32'h00000000;
    weight_mem[1135] = 32'h00000000;
    weight_mem[1136] = 32'h00000000;
    weight_mem[1137] = 32'h00000000;
    weight_mem[1138] = 32'h00000000;
    weight_mem[1139] = 32'h00000000;
    weight_mem[1140] = 32'h00000000;
    weight_mem[1141] = 32'h00000000;
    weight_mem[1142] = 32'h00000000;
    weight_mem[1143] = 32'h00000000;
    weight_mem[1144] = 32'h00000000;
    weight_mem[1145] = 32'h00000000;
    weight_mem[1146] = 32'h00000000;
    weight_mem[1147] = 32'h00000000;
    weight_mem[1148] = 32'h00000000;
    weight_mem[1149] = 32'h00000000;
    weight_mem[1150] = 32'h00000000;
    weight_mem[1151] = 32'h00000000;
    weight_mem[1152] = 32'h00000000;
    weight_mem[1153] = 32'h00000000;
    weight_mem[1154] = 32'h00000000;
    weight_mem[1155] = 32'h00000000;
    weight_mem[1156] = 32'h00000000;
    weight_mem[1157] = 32'h00000000;
    weight_mem[1158] = 32'h00000000;
    weight_mem[1159] = 32'h00000000;
    weight_mem[1160] = 32'h00000000;
    weight_mem[1161] = 32'h00000000;
    weight_mem[1162] = 32'h00000000;
    weight_mem[1163] = 32'h00000000;
    weight_mem[1164] = 32'h00000000;
    weight_mem[1165] = 32'h00000000;
    weight_mem[1166] = 32'h00000000;
    weight_mem[1167] = 32'h00000000;
    weight_mem[1168] = 32'h00000000;
    weight_mem[1169] = 32'h00000000;
    weight_mem[1170] = 32'h00000000;
    weight_mem[1171] = 32'h00000000;
    weight_mem[1172] = 32'h00000000;
    weight_mem[1173] = 32'h00000000;
    weight_mem[1174] = 32'h00000000;
    weight_mem[1175] = 32'h00000000;
    weight_mem[1176] = 32'h00000000;
    weight_mem[1177] = 32'h00000000;
    weight_mem[1178] = 32'h00000000;
    weight_mem[1179] = 32'h00000000;
    weight_mem[1180] = 32'h00000000;
    weight_mem[1181] = 32'h00000000;
    weight_mem[1182] = 32'h00000000;
    weight_mem[1183] = 32'h00000000;
    weight_mem[1184] = 32'h00000000;
    weight_mem[1185] = 32'h00000000;
    weight_mem[1186] = 32'h00000000;
    weight_mem[1187] = 32'h00000000;
    weight_mem[1188] = 32'h00000000;
    weight_mem[1189] = 32'h00000000;
    weight_mem[1190] = 32'h00000000;
    weight_mem[1191] = 32'h00000000;
    weight_mem[1192] = 32'h00000000;
    weight_mem[1193] = 32'h00000000;
    weight_mem[1194] = 32'h00000000;
    weight_mem[1195] = 32'h00000000;
    weight_mem[1196] = 32'h00000000;
    weight_mem[1197] = 32'h00000000;
    weight_mem[1198] = 32'h00000000;
    weight_mem[1199] = 32'h00000000;
    weight_mem[1200] = 32'h00000000;
    weight_mem[1201] = 32'h00000000;
    weight_mem[1202] = 32'h00000000;
    weight_mem[1203] = 32'h00000000;
    weight_mem[1204] = 32'h00000000;
    weight_mem[1205] = 32'h00000000;
    weight_mem[1206] = 32'h00000000;
    weight_mem[1207] = 32'h00000000;
    weight_mem[1208] = 32'h00000000;
    weight_mem[1209] = 32'h00000000;
    weight_mem[1210] = 32'h00000000;
    weight_mem[1211] = 32'h00000000;
    weight_mem[1212] = 32'h00000000;
    weight_mem[1213] = 32'h00000000;
    weight_mem[1214] = 32'h00000000;
    weight_mem[1215] = 32'h00000000;
    weight_mem[1216] = 32'h00000000;
    weight_mem[1217] = 32'h00000000;
    weight_mem[1218] = 32'h00000000;
    weight_mem[1219] = 32'h00000000;
    weight_mem[1220] = 32'h00000000;
    weight_mem[1221] = 32'h00000000;
    weight_mem[1222] = 32'h00000000;
    weight_mem[1223] = 32'h00000000;
    weight_mem[1224] = 32'h00000000;
    weight_mem[1225] = 32'h00000000;
    weight_mem[1226] = 32'h00000000;
    weight_mem[1227] = 32'h00000000;
    weight_mem[1228] = 32'h00000000;
    weight_mem[1229] = 32'h00000000;
    weight_mem[1230] = 32'h00000000;
    weight_mem[1231] = 32'h00000000;
    weight_mem[1232] = 32'h00000000;
    weight_mem[1233] = 32'h00000000;
    weight_mem[1234] = 32'h00000000;
    weight_mem[1235] = 32'h00000000;
    weight_mem[1236] = 32'h00000000;
    weight_mem[1237] = 32'h00000000;
    weight_mem[1238] = 32'h00000000;
    weight_mem[1239] = 32'h00000000;
    weight_mem[1240] = 32'h00000000;
    weight_mem[1241] = 32'h00000000;
    weight_mem[1242] = 32'h00000000;
    weight_mem[1243] = 32'h00000000;
    weight_mem[1244] = 32'h00000000;
    weight_mem[1245] = 32'h00000000;
    weight_mem[1246] = 32'h00000000;
    weight_mem[1247] = 32'h00000000;
    weight_mem[1248] = 32'h00000000;
    weight_mem[1249] = 32'h00000000;
    weight_mem[1250] = 32'h00000000;
    weight_mem[1251] = 32'h00000000;
    weight_mem[1252] = 32'h00000000;
    weight_mem[1253] = 32'h00000000;
    weight_mem[1254] = 32'h00000000;
    weight_mem[1255] = 32'h00000000;
    weight_mem[1256] = 32'h00000000;
    weight_mem[1257] = 32'h00000000;
    weight_mem[1258] = 32'h00000000;
    weight_mem[1259] = 32'h00000000;
    weight_mem[1260] = 32'h00000000;
    weight_mem[1261] = 32'h00000000;
    weight_mem[1262] = 32'h00000000;
    weight_mem[1263] = 32'h00000000;
    weight_mem[1264] = 32'h00000000;
    weight_mem[1265] = 32'h00000000;
    weight_mem[1266] = 32'h00000000;
    weight_mem[1267] = 32'h00000000;
    weight_mem[1268] = 32'h00000000;
    weight_mem[1269] = 32'h00000000;
    weight_mem[1270] = 32'h00000000;
    weight_mem[1271] = 32'h00000000;
    weight_mem[1272] = 32'h00000000;
    weight_mem[1273] = 32'h00000000;
    weight_mem[1274] = 32'h00000000;
    weight_mem[1275] = 32'h00000000;
    weight_mem[1276] = 32'h00000000;
    weight_mem[1277] = 32'h00000000;
    weight_mem[1278] = 32'h00000000;
    weight_mem[1279] = 32'h00000000;
    weight_mem[1280] = 32'h00000000;
    weight_mem[1281] = 32'h00000000;
    weight_mem[1282] = 32'h00000000;
end

initial begin
    weight_b_mem[0] = 32'h00000000;
    weight_b_mem[1] = 32'h00000000;
    weight_b_mem[2] = 32'h00000000;
    weight_b_mem[3] = 32'h00000000;
    weight_b_mem[4] = 32'h00000000;
    weight_b_mem[5] = 32'h00000000;
    weight_b_mem[6] = 32'h00000000;
    weight_b_mem[7] = 32'h00000000;
    weight_b_mem[8] = 32'h00000000;
    weight_b_mem[9] = 32'h00000000;
    weight_b_mem[10] = 32'h00000000;
    weight_b_mem[11] = 32'h00000000;
    weight_b_mem[12] = 32'h00000000;
    weight_b_mem[13] = 32'h00000000;
    weight_b_mem[14] = 32'h00000000;
    weight_b_mem[15] = 32'h00000000;
    weight_b_mem[16] = 32'h00000000;
    weight_b_mem[17] = 32'h00000000;
    weight_b_mem[18] = 32'h00000000;
    weight_b_mem[19] = 32'h00000000;
    weight_b_mem[20] = 32'h00000000;
    weight_b_mem[21] = 32'h00000000;
    weight_b_mem[22] = 32'h00000000;
    weight_b_mem[23] = 32'h00000000;
    weight_b_mem[24] = 32'h00000000;
    weight_b_mem[25] = 32'h00000000;
    weight_b_mem[26] = 32'h00000000;
    weight_b_mem[27] = 32'h00000000;
    weight_b_mem[28] = 32'h00000000;
    weight_b_mem[29] = 32'h00000000;
    weight_b_mem[30] = 32'h00000000;
    weight_b_mem[31] = 32'h00000000;
    weight_b_mem[32] = 32'h00000000;
    weight_b_mem[33] = 32'h00000000;
    weight_b_mem[34] = 32'h00000000;
    weight_b_mem[35] = 32'h00000000;
    weight_b_mem[36] = 32'h00000000;
    weight_b_mem[37] = 32'h00000000;
    weight_b_mem[38] = 32'h00000000;
    weight_b_mem[39] = 32'h00000000;
    weight_b_mem[40] = 32'h00000000;
    weight_b_mem[41] = 32'h00000000;
    weight_b_mem[42] = 32'h00000000;
    weight_b_mem[43] = 32'h00000000;
    weight_b_mem[44] = 32'h00000000;
    weight_b_mem[45] = 32'h00000000;
    weight_b_mem[46] = 32'h00000000;
    weight_b_mem[47] = 32'h00000000;
    weight_b_mem[48] = 32'h00000000;
    weight_b_mem[49] = 32'h00000000;
    weight_b_mem[50] = 32'h00000000;
    weight_b_mem[51] = 32'h00000000;
    weight_b_mem[52] = 32'h00000000;
    weight_b_mem[53] = 32'h00000000;
    weight_b_mem[54] = 32'h00000000;
    weight_b_mem[55] = 32'h00000000;
    weight_b_mem[56] = 32'h00000000;
    weight_b_mem[57] = 32'h00000000;
    weight_b_mem[58] = 32'h00000000;
    weight_b_mem[59] = 32'h00000000;
    weight_b_mem[60] = 32'h00000000;
    weight_b_mem[61] = 32'h00000000;
    weight_b_mem[62] = 32'h00000000;
    weight_b_mem[63] = 32'h00000000;
    weight_b_mem[64] = 32'h00000000;
    weight_b_mem[65] = 32'h00000000;
    weight_b_mem[66] = 32'h00000000;
    weight_b_mem[67] = 32'h00000000;
    weight_b_mem[68] = 32'h00000000;
    weight_b_mem[69] = 32'h00000000;
    weight_b_mem[70] = 32'h00000000;
    weight_b_mem[71] = 32'h00000000;
    weight_b_mem[72] = 32'h00000000;
    weight_b_mem[73] = 32'h00000000;
    weight_b_mem[74] = 32'h00000000;
    weight_b_mem[75] = 32'h00000000;
    weight_b_mem[76] = 32'h00000000;
    weight_b_mem[77] = 32'h00000000;
    weight_b_mem[78] = 32'h00000000;
    weight_b_mem[79] = 32'h00000000;
    weight_b_mem[80] = 32'h00000000;
    weight_b_mem[81] = 32'h00000000;
    weight_b_mem[82] = 32'h00000000;
    weight_b_mem[83] = 32'h00000000;
    weight_b_mem[84] = 32'h00000000;
    weight_b_mem[85] = 32'h00000000;
    weight_b_mem[86] = 32'h00000000;
    weight_b_mem[87] = 32'h00000000;
    weight_b_mem[88] = 32'h00000000;
    weight_b_mem[89] = 32'h00000000;
    weight_b_mem[90] = 32'h00000000;
    weight_b_mem[91] = 32'h00000000;
    weight_b_mem[92] = 32'h00000000;
    weight_b_mem[93] = 32'h00000000;
    weight_b_mem[94] = 32'h00000000;
    weight_b_mem[95] = 32'h00000000;
    weight_b_mem[96] = 32'h00000000;
    weight_b_mem[97] = 32'h00000000;
    weight_b_mem[98] = 32'h00000000;
    weight_b_mem[99] = 32'h00000000;
    weight_b_mem[100] = 32'h00000000;
    weight_b_mem[101] = 32'h00000000;
    weight_b_mem[102] = 32'h00000000;
    weight_b_mem[103] = 32'h00000000;
    weight_b_mem[104] = 32'h00000000;
    weight_b_mem[105] = 32'h00000000;
    weight_b_mem[106] = 32'h00000000;
    weight_b_mem[107] = 32'h00000000;
    weight_b_mem[108] = 32'h00000000;
    weight_b_mem[109] = 32'h00000000;
    weight_b_mem[110] = 32'h00000000;
    weight_b_mem[111] = 32'h00000000;
    weight_b_mem[112] = 32'h00000000;
    weight_b_mem[113] = 32'h00000000;
    weight_b_mem[114] = 32'h00000000;
    weight_b_mem[115] = 32'h00000000;
    weight_b_mem[116] = 32'h00000000;
    weight_b_mem[117] = 32'h00000000;
    weight_b_mem[118] = 32'h00000000;
    weight_b_mem[119] = 32'h00000000;
    weight_b_mem[120] = 32'h00000000;
    weight_b_mem[121] = 32'h00000000;
    weight_b_mem[122] = 32'h00000000;
    weight_b_mem[123] = 32'h00000000;
    weight_b_mem[124] = 32'h00000000;
    weight_b_mem[125] = 32'h00000000;
    weight_b_mem[126] = 32'h00000000;
    weight_b_mem[127] = 32'h00000000;
    weight_b_mem[128] = 32'h00000000;
    weight_b_mem[129] = 32'h00000000;
    weight_b_mem[130] = 32'h00000000;
    weight_b_mem[131] = 32'h00000000;
    weight_b_mem[132] = 32'h00000000;
    weight_b_mem[133] = 32'h00000000;
    weight_b_mem[134] = 32'h00000000;
    weight_b_mem[135] = 32'h00000000;
    weight_b_mem[136] = 32'h00000000;
    weight_b_mem[137] = 32'h00000000;
    weight_b_mem[138] = 32'h00000000;
    weight_b_mem[139] = 32'h00000000;
    weight_b_mem[140] = 32'h00000000;
    weight_b_mem[141] = 32'h00000000;
    weight_b_mem[142] = 32'h00000000;
    weight_b_mem[143] = 32'h00000000;
    weight_b_mem[144] = 32'h00000000;
    weight_b_mem[145] = 32'h00000000;
    weight_b_mem[146] = 32'h00000000;
    weight_b_mem[147] = 32'h00000000;
    weight_b_mem[148] = 32'h00000000;
    weight_b_mem[149] = 32'h00000000;
    weight_b_mem[150] = 32'h00000000;
    weight_b_mem[151] = 32'h00000000;
    weight_b_mem[152] = 32'h00000000;
    weight_b_mem[153] = 32'h00000000;
    weight_b_mem[154] = 32'h00000000;
    weight_b_mem[155] = 32'h00000000;
    weight_b_mem[156] = 32'h00000000;
    weight_b_mem[157] = 32'h00000000;
    weight_b_mem[158] = 32'h00000000;
    weight_b_mem[159] = 32'h00000000;
    weight_b_mem[160] = 32'h00000000;
    weight_b_mem[161] = 32'h00000000;
    weight_b_mem[162] = 32'h00000000;
    weight_b_mem[163] = 32'h00000000;
    weight_b_mem[164] = 32'h00000000;
    weight_b_mem[165] = 32'h00000000;
    weight_b_mem[166] = 32'h00000000;
    weight_b_mem[167] = 32'h00000000;
    weight_b_mem[168] = 32'h00000000;
    weight_b_mem[169] = 32'h00000000;
    weight_b_mem[170] = 32'h00000000;
    weight_b_mem[171] = 32'h00000000;
    weight_b_mem[172] = 32'h00000000;
    weight_b_mem[173] = 32'h00000000;
    weight_b_mem[174] = 32'h00000000;
    weight_b_mem[175] = 32'h00000000;
    weight_b_mem[176] = 32'h00000000;
    weight_b_mem[177] = 32'h00000000;
    weight_b_mem[178] = 32'h00000000;
    weight_b_mem[179] = 32'h00000000;
    weight_b_mem[180] = 32'h00000000;
    weight_b_mem[181] = 32'h00000000;
    weight_b_mem[182] = 32'h00000000;
    weight_b_mem[183] = 32'h00000000;
    weight_b_mem[184] = 32'h00000000;
    weight_b_mem[185] = 32'h00000000;
    weight_b_mem[186] = 32'h00000000;
    weight_b_mem[187] = 32'h00000000;
    weight_b_mem[188] = 32'h00000000;
    weight_b_mem[189] = 32'h00000000;
    weight_b_mem[190] = 32'h00000000;
    weight_b_mem[191] = 32'h00000000;
    weight_b_mem[192] = 32'h00000000;
    weight_b_mem[193] = 32'h00000000;
    weight_b_mem[194] = 32'h00000000;
    weight_b_mem[195] = 32'h00000000;
    weight_b_mem[196] = 32'h00000000;
    weight_b_mem[197] = 32'h00000000;
    weight_b_mem[198] = 32'h00000000;
    weight_b_mem[199] = 32'h00000000;
    weight_b_mem[200] = 32'h00000000;
    weight_b_mem[201] = 32'h00000000;
    weight_b_mem[202] = 32'h00000000;
    weight_b_mem[203] = 32'h00000000;
    weight_b_mem[204] = 32'h00000000;
    weight_b_mem[205] = 32'h00000000;
    weight_b_mem[206] = 32'h00000000;
    weight_b_mem[207] = 32'h00000000;
    weight_b_mem[208] = 32'h00000000;
    weight_b_mem[209] = 32'h00000000;
    weight_b_mem[210] = 32'h00000000;
    weight_b_mem[211] = 32'h00000000;
    weight_b_mem[212] = 32'h00000000;
    weight_b_mem[213] = 32'h00000000;
    weight_b_mem[214] = 32'h00000000;
    weight_b_mem[215] = 32'h00000000;
    weight_b_mem[216] = 32'h00000000;
    weight_b_mem[217] = 32'h00000000;
    weight_b_mem[218] = 32'h00000000;
    weight_b_mem[219] = 32'h00000000;
    weight_b_mem[220] = 32'h00000000;
    weight_b_mem[221] = 32'h00000000;
    weight_b_mem[222] = 32'h00000000;
    weight_b_mem[223] = 32'h00000000;
    weight_b_mem[224] = 32'h00000000;
    weight_b_mem[225] = 32'h00000000;
    weight_b_mem[226] = 32'h00000000;
    weight_b_mem[227] = 32'h00000000;
    weight_b_mem[228] = 32'h00000000;
    weight_b_mem[229] = 32'h00000000;
    weight_b_mem[230] = 32'h00000000;
    weight_b_mem[231] = 32'h00000000;
    weight_b_mem[232] = 32'h00000000;
    weight_b_mem[233] = 32'h00000000;
    weight_b_mem[234] = 32'h00000000;
    weight_b_mem[235] = 32'h00000000;
    weight_b_mem[236] = 32'h00000000;
    weight_b_mem[237] = 32'h00000000;
    weight_b_mem[238] = 32'h00000000;
    weight_b_mem[239] = 32'h00000000;
    weight_b_mem[240] = 32'h00000000;
    weight_b_mem[241] = 32'h00000000;
    weight_b_mem[242] = 32'h00000000;
    weight_b_mem[243] = 32'h00000000;
    weight_b_mem[244] = 32'h00000000;
    weight_b_mem[245] = 32'h00000000;
    weight_b_mem[246] = 32'h00000000;
    weight_b_mem[247] = 32'h00000000;
    weight_b_mem[248] = 32'h00000000;
    weight_b_mem[249] = 32'h00000000;
    weight_b_mem[250] = 32'h00000000;
    weight_b_mem[251] = 32'h00000000;
    weight_b_mem[252] = 32'h00000000;
    weight_b_mem[253] = 32'h00000000;
    weight_b_mem[254] = 32'h00000000;
    weight_b_mem[255] = 32'h00000000;
    weight_b_mem[256] = 32'h00000000;
    weight_b_mem[257] = 32'h00000000;
    weight_b_mem[258] = 32'h00000000;
    weight_b_mem[259] = 32'h00000000;
    weight_b_mem[260] = 32'h00000000;
    weight_b_mem[261] = 32'h00000000;
    weight_b_mem[262] = 32'h00000000;
    weight_b_mem[263] = 32'h00000000;
    weight_b_mem[264] = 32'h00000000;
    weight_b_mem[265] = 32'h00000000;
    weight_b_mem[266] = 32'h00000000;
    weight_b_mem[267] = 32'h00000000;
    weight_b_mem[268] = 32'h00000000;
    weight_b_mem[269] = 32'h00000000;
    weight_b_mem[270] = 32'h00000000;
    weight_b_mem[271] = 32'h00000000;
    weight_b_mem[272] = 32'h00000000;
    weight_b_mem[273] = 32'h00000000;
    weight_b_mem[274] = 32'h00000000;
    weight_b_mem[275] = 32'h00000000;
    weight_b_mem[276] = 32'h00000000;
    weight_b_mem[277] = 32'h00000000;
    weight_b_mem[278] = 32'h00000000;
    weight_b_mem[279] = 32'h00000000;
    weight_b_mem[280] = 32'h00000000;
    weight_b_mem[281] = 32'h00000000;
    weight_b_mem[282] = 32'h00000000;
    weight_b_mem[283] = 32'h00000000;
    weight_b_mem[284] = 32'h00000000;
    weight_b_mem[285] = 32'h00000000;
    weight_b_mem[286] = 32'h00000000;
    weight_b_mem[287] = 32'h00000000;
    weight_b_mem[288] = 32'h00000000;
    weight_b_mem[289] = 32'h00000000;
    weight_b_mem[290] = 32'h00000000;
    weight_b_mem[291] = 32'h00000000;
    weight_b_mem[292] = 32'h00000000;
    weight_b_mem[293] = 32'h00000000;
    weight_b_mem[294] = 32'h00000000;
    weight_b_mem[295] = 32'h00000000;
    weight_b_mem[296] = 32'h00000000;
    weight_b_mem[297] = 32'h00000000;
    weight_b_mem[298] = 32'h00000000;
    weight_b_mem[299] = 32'h00000000;
    weight_b_mem[300] = 32'h00000000;
    weight_b_mem[301] = 32'h00000000;
    weight_b_mem[302] = 32'h00000000;
    weight_b_mem[303] = 32'h00000000;
    weight_b_mem[304] = 32'h00000000;
    weight_b_mem[305] = 32'h00000000;
    weight_b_mem[306] = 32'h00000000;
    weight_b_mem[307] = 32'h00000000;
    weight_b_mem[308] = 32'h00000000;
    weight_b_mem[309] = 32'h00000000;
    weight_b_mem[310] = 32'h00000000;
    weight_b_mem[311] = 32'h00000000;
    weight_b_mem[312] = 32'h00000000;
    weight_b_mem[313] = 32'h00000000;
    weight_b_mem[314] = 32'h00000000;
    weight_b_mem[315] = 32'h00000000;
    weight_b_mem[316] = 32'h00000000;
    weight_b_mem[317] = 32'h00000000;
    weight_b_mem[318] = 32'h00000000;
    weight_b_mem[319] = 32'h00000000;
    weight_b_mem[320] = 32'h00000000;
    weight_b_mem[321] = 32'h00000000;
    weight_b_mem[322] = 32'h00000000;
    weight_b_mem[323] = 32'h00000000;
    weight_b_mem[324] = 32'h00000000;
    weight_b_mem[325] = 32'h00000000;
    weight_b_mem[326] = 32'h00000000;
    weight_b_mem[327] = 32'h00000000;
    weight_b_mem[328] = 32'h00000000;
    weight_b_mem[329] = 32'h00000000;
    weight_b_mem[330] = 32'h00000000;
    weight_b_mem[331] = 32'h00000000;
    weight_b_mem[332] = 32'h00000000;
    weight_b_mem[333] = 32'h00000000;
    weight_b_mem[334] = 32'h00000000;
    weight_b_mem[335] = 32'h00000000;
    weight_b_mem[336] = 32'h00000000;
    weight_b_mem[337] = 32'h00000000;
    weight_b_mem[338] = 32'h00000000;
    weight_b_mem[339] = 32'h00000000;
    weight_b_mem[340] = 32'h00000000;
    weight_b_mem[341] = 32'h00000000;
    weight_b_mem[342] = 32'h00000000;
    weight_b_mem[343] = 32'h00000000;
    weight_b_mem[344] = 32'h00000000;
    weight_b_mem[345] = 32'h00000000;
    weight_b_mem[346] = 32'h00000000;
    weight_b_mem[347] = 32'h00000000;
    weight_b_mem[348] = 32'h00000000;
    weight_b_mem[349] = 32'h00000000;
    weight_b_mem[350] = 32'h00000000;
    weight_b_mem[351] = 32'h00000000;
    weight_b_mem[352] = 32'h00000000;
    weight_b_mem[353] = 32'h00000000;
    weight_b_mem[354] = 32'h00000000;
    weight_b_mem[355] = 32'h00000000;
    weight_b_mem[356] = 32'h00000000;
    weight_b_mem[357] = 32'h00000000;
    weight_b_mem[358] = 32'h00000000;
    weight_b_mem[359] = 32'h00000000;
    weight_b_mem[360] = 32'h00000000;
    weight_b_mem[361] = 32'h00000000;
    weight_b_mem[362] = 32'h00000000;
    weight_b_mem[363] = 32'h00000000;
    weight_b_mem[364] = 32'h00000000;
    weight_b_mem[365] = 32'h00000000;
    weight_b_mem[366] = 32'h00000000;
    weight_b_mem[367] = 32'h00000000;
    weight_b_mem[368] = 32'h00000000;
    weight_b_mem[369] = 32'h00000000;
    weight_b_mem[370] = 32'h00000000;
    weight_b_mem[371] = 32'h00000000;
    weight_b_mem[372] = 32'h00000000;
    weight_b_mem[373] = 32'h00000000;
    weight_b_mem[374] = 32'h00000000;
    weight_b_mem[375] = 32'h00000000;
    weight_b_mem[376] = 32'h00000000;
    weight_b_mem[377] = 32'h00000000;
    weight_b_mem[378] = 32'h00000000;
    weight_b_mem[379] = 32'h00000000;
    weight_b_mem[380] = 32'h00000000;
    weight_b_mem[381] = 32'h00000000;
    weight_b_mem[382] = 32'h00000000;
    weight_b_mem[383] = 32'h00000000;
    weight_b_mem[384] = 32'h00000000;
    weight_b_mem[385] = 32'h00000000;
    weight_b_mem[386] = 32'h00000000;
    weight_b_mem[387] = 32'h00000000;
    weight_b_mem[388] = 32'h00000000;
    weight_b_mem[389] = 32'h00000000;
    weight_b_mem[390] = 32'h00000000;
    weight_b_mem[391] = 32'h00000000;
    weight_b_mem[392] = 32'h00000000;
    weight_b_mem[393] = 32'h00000000;
    weight_b_mem[394] = 32'h00000000;
    weight_b_mem[395] = 32'h00000000;
    weight_b_mem[396] = 32'h00000000;
    weight_b_mem[397] = 32'h00000000;
    weight_b_mem[398] = 32'h00000000;
    weight_b_mem[399] = 32'h00000000;
    weight_b_mem[400] = 32'h00000000;
    weight_b_mem[401] = 32'h00000000;
    weight_b_mem[402] = 32'h00000000;
    weight_b_mem[403] = 32'h00000000;
    weight_b_mem[404] = 32'h00000000;
    weight_b_mem[405] = 32'h00000000;
    weight_b_mem[406] = 32'h00000000;
    weight_b_mem[407] = 32'h00000000;
    weight_b_mem[408] = 32'h00000000;
    weight_b_mem[409] = 32'h00000000;
    weight_b_mem[410] = 32'h00000000;
    weight_b_mem[411] = 32'h00000000;
    weight_b_mem[412] = 32'h00000000;
    weight_b_mem[413] = 32'h00000000;
    weight_b_mem[414] = 32'h00000000;
    weight_b_mem[415] = 32'h00000000;
    weight_b_mem[416] = 32'h00000000;
    weight_b_mem[417] = 32'h00000000;
    weight_b_mem[418] = 32'h00000000;
    weight_b_mem[419] = 32'h00000000;
    weight_b_mem[420] = 32'h00000000;
    weight_b_mem[421] = 32'h00000000;
    weight_b_mem[422] = 32'h00000000;
    weight_b_mem[423] = 32'h00000000;
    weight_b_mem[424] = 32'h00000000;
    weight_b_mem[425] = 32'h00000000;
    weight_b_mem[426] = 32'h00000000;
    weight_b_mem[427] = 32'h00000000;
    weight_b_mem[428] = 32'h00000000;
    weight_b_mem[429] = 32'h00000000;
    weight_b_mem[430] = 32'h00000000;
    weight_b_mem[431] = 32'h00000000;
    weight_b_mem[432] = 32'h00000000;
    weight_b_mem[433] = 32'h00000000;
    weight_b_mem[434] = 32'h00000000;
    weight_b_mem[435] = 32'h00000000;
    weight_b_mem[436] = 32'h00000000;
    weight_b_mem[437] = 32'h00000000;
    weight_b_mem[438] = 32'h00000000;
    weight_b_mem[439] = 32'h00000000;
    weight_b_mem[440] = 32'h00000000;
    weight_b_mem[441] = 32'h00000000;
    weight_b_mem[442] = 32'h00000000;
    weight_b_mem[443] = 32'h00000000;
    weight_b_mem[444] = 32'h00000000;
    weight_b_mem[445] = 32'h00000000;
    weight_b_mem[446] = 32'h00000000;
    weight_b_mem[447] = 32'h00000000;
    weight_b_mem[448] = 32'h00000000;
    weight_b_mem[449] = 32'h00000000;
    weight_b_mem[450] = 32'h00000000;
    weight_b_mem[451] = 32'h00000000;
    weight_b_mem[452] = 32'h00000000;
    weight_b_mem[453] = 32'h00000000;
    weight_b_mem[454] = 32'h00000000;
    weight_b_mem[455] = 32'h00000000;
    weight_b_mem[456] = 32'h00000000;
    weight_b_mem[457] = 32'h00000000;
    weight_b_mem[458] = 32'h00000000;
    weight_b_mem[459] = 32'h00000000;
    weight_b_mem[460] = 32'h00000000;
    weight_b_mem[461] = 32'h00000000;
    weight_b_mem[462] = 32'h00000000;
    weight_b_mem[463] = 32'h00000000;
    weight_b_mem[464] = 32'h00000000;
    weight_b_mem[465] = 32'h00000000;
    weight_b_mem[466] = 32'h00000000;
    weight_b_mem[467] = 32'h00000000;
    weight_b_mem[468] = 32'h00000000;
    weight_b_mem[469] = 32'h00000000;
    weight_b_mem[470] = 32'h00000000;
    weight_b_mem[471] = 32'h00000000;
    weight_b_mem[472] = 32'h00000000;
    weight_b_mem[473] = 32'h00000000;
    weight_b_mem[474] = 32'h00000000;
    weight_b_mem[475] = 32'h00000000;
    weight_b_mem[476] = 32'h00000000;
    weight_b_mem[477] = 32'h00000000;
    weight_b_mem[478] = 32'h00000000;
    weight_b_mem[479] = 32'h00000000;
    weight_b_mem[480] = 32'h00000000;
    weight_b_mem[481] = 32'h00000000;
    weight_b_mem[482] = 32'h00000000;
    weight_b_mem[483] = 32'h00000000;
    weight_b_mem[484] = 32'h00000000;
    weight_b_mem[485] = 32'h00000000;
    weight_b_mem[486] = 32'h00000000;
    weight_b_mem[487] = 32'h00000000;
    weight_b_mem[488] = 32'h00000000;
    weight_b_mem[489] = 32'h00000000;
    weight_b_mem[490] = 32'h00000000;
    weight_b_mem[491] = 32'h00000000;
    weight_b_mem[492] = 32'h00000000;
    weight_b_mem[493] = 32'h00000000;
    weight_b_mem[494] = 32'h00000000;
    weight_b_mem[495] = 32'h00000000;
    weight_b_mem[496] = 32'h00000000;
    weight_b_mem[497] = 32'h00000000;
    weight_b_mem[498] = 32'h00000000;
    weight_b_mem[499] = 32'h00000000;
    weight_b_mem[500] = 32'h00000000;
    weight_b_mem[501] = 32'h00000000;
    weight_b_mem[502] = 32'h00000000;
    weight_b_mem[503] = 32'h00000000;
    weight_b_mem[504] = 32'h00000000;
    weight_b_mem[505] = 32'h00000000;
    weight_b_mem[506] = 32'h00000000;
    weight_b_mem[507] = 32'h00000000;
    weight_b_mem[508] = 32'h00000000;
    weight_b_mem[509] = 32'h00000000;
    weight_b_mem[510] = 32'h00000000;
    weight_b_mem[511] = 32'h00000000;
    weight_b_mem[512] = 32'h00000000;
    weight_b_mem[513] = 32'h00000000;
    weight_b_mem[514] = 32'h00000000;
    weight_b_mem[515] = 32'h00000000;
    weight_b_mem[516] = 32'h00000000;
    weight_b_mem[517] = 32'h00000000;
    weight_b_mem[518] = 32'h00000000;
    weight_b_mem[519] = 32'h00000000;
    weight_b_mem[520] = 32'h00000000;
    weight_b_mem[521] = 32'h00000000;
    weight_b_mem[522] = 32'h00000000;
    weight_b_mem[523] = 32'h00000000;
    weight_b_mem[524] = 32'h00000000;
    weight_b_mem[525] = 32'h00000000;
    weight_b_mem[526] = 32'h00000000;
    weight_b_mem[527] = 32'h00000000;
    weight_b_mem[528] = 32'h00000000;
    weight_b_mem[529] = 32'h00000000;
    weight_b_mem[530] = 32'h00000000;
    weight_b_mem[531] = 32'h00000000;
    weight_b_mem[532] = 32'h00000000;
    weight_b_mem[533] = 32'h00000000;
    weight_b_mem[534] = 32'h00000000;
    weight_b_mem[535] = 32'h00000000;
    weight_b_mem[536] = 32'h00000000;
    weight_b_mem[537] = 32'h00000000;
    weight_b_mem[538] = 32'h00000000;
    weight_b_mem[539] = 32'h00000000;
    weight_b_mem[540] = 32'h00000000;
    weight_b_mem[541] = 32'h00000000;
    weight_b_mem[542] = 32'h00000000;
    weight_b_mem[543] = 32'h00000000;
    weight_b_mem[544] = 32'h00000000;
    weight_b_mem[545] = 32'h00000000;
    weight_b_mem[546] = 32'h00000000;
    weight_b_mem[547] = 32'h00000000;
    weight_b_mem[548] = 32'h00000000;
    weight_b_mem[549] = 32'h00000000;
    weight_b_mem[550] = 32'h00000000;
    weight_b_mem[551] = 32'h00000000;
    weight_b_mem[552] = 32'h00000000;
    weight_b_mem[553] = 32'h00000000;
    weight_b_mem[554] = 32'h00000000;
    weight_b_mem[555] = 32'h00000000;
    weight_b_mem[556] = 32'h00000000;
    weight_b_mem[557] = 32'h00000000;
    weight_b_mem[558] = 32'h00000000;
    weight_b_mem[559] = 32'h00000000;
    weight_b_mem[560] = 32'h00000000;
    weight_b_mem[561] = 32'h00000000;
    weight_b_mem[562] = 32'h00000000;
    weight_b_mem[563] = 32'h00000000;
    weight_b_mem[564] = 32'h00000000;
    weight_b_mem[565] = 32'h00000000;
    weight_b_mem[566] = 32'h00000000;
    weight_b_mem[567] = 32'h00000000;
    weight_b_mem[568] = 32'h00000000;
    weight_b_mem[569] = 32'h00000000;
    weight_b_mem[570] = 32'h00000000;
    weight_b_mem[571] = 32'h00000000;
    weight_b_mem[572] = 32'h00000000;
    weight_b_mem[573] = 32'h00000000;
    weight_b_mem[574] = 32'h00000000;
    weight_b_mem[575] = 32'h00000000;
    weight_b_mem[576] = 32'h00000000;
    weight_b_mem[577] = 32'h00000000;
    weight_b_mem[578] = 32'h00000000;
    weight_b_mem[579] = 32'h00000000;
    weight_b_mem[580] = 32'h00000000;
    weight_b_mem[581] = 32'h00000000;
    weight_b_mem[582] = 32'h00000000;
    weight_b_mem[583] = 32'h00000000;
    weight_b_mem[584] = 32'h00000000;
    weight_b_mem[585] = 32'h00000000;
    weight_b_mem[586] = 32'h00000000;
    weight_b_mem[587] = 32'h00000000;
    weight_b_mem[588] = 32'h00000000;
    weight_b_mem[589] = 32'h00000000;
    weight_b_mem[590] = 32'h00000000;
    weight_b_mem[591] = 32'h00000000;
    weight_b_mem[592] = 32'h00000000;
    weight_b_mem[593] = 32'h00000000;
    weight_b_mem[594] = 32'h00000000;
    weight_b_mem[595] = 32'h00000000;
    weight_b_mem[596] = 32'h00000000;
    weight_b_mem[597] = 32'h00000000;
    weight_b_mem[598] = 32'h00000000;
    weight_b_mem[599] = 32'h00000000;
    weight_b_mem[600] = 32'h00000000;
    weight_b_mem[601] = 32'h00000000;
    weight_b_mem[602] = 32'h00000000;
    weight_b_mem[603] = 32'h00000000;
    weight_b_mem[604] = 32'h00000000;
    weight_b_mem[605] = 32'h00000000;
    weight_b_mem[606] = 32'h00000000;
    weight_b_mem[607] = 32'h00000000;
    weight_b_mem[608] = 32'h00000000;
    weight_b_mem[609] = 32'h00000000;
    weight_b_mem[610] = 32'h00000000;
    weight_b_mem[611] = 32'h00000000;
    weight_b_mem[612] = 32'h00000000;
    weight_b_mem[613] = 32'h00000000;
    weight_b_mem[614] = 32'h00000000;
    weight_b_mem[615] = 32'h00000000;
    weight_b_mem[616] = 32'h00000000;
    weight_b_mem[617] = 32'h00000000;
    weight_b_mem[618] = 32'h00000000;
    weight_b_mem[619] = 32'h00000000;
    weight_b_mem[620] = 32'h00000000;
    weight_b_mem[621] = 32'h00000000;
    weight_b_mem[622] = 32'h00000000;
    weight_b_mem[623] = 32'h00000000;
    weight_b_mem[624] = 32'h00000000;
    weight_b_mem[625] = 32'h00000000;
    weight_b_mem[626] = 32'h00000000;
    weight_b_mem[627] = 32'h00000000;
    weight_b_mem[628] = 32'h00000000;
    weight_b_mem[629] = 32'h00000000;
    weight_b_mem[630] = 32'h00000000;
    weight_b_mem[631] = 32'h00000000;
    weight_b_mem[632] = 32'h00000000;
    weight_b_mem[633] = 32'h00000000;
    weight_b_mem[634] = 32'h00000000;
    weight_b_mem[635] = 32'h00000000;
    weight_b_mem[636] = 32'h00000000;
    weight_b_mem[637] = 32'h00000000;
    weight_b_mem[638] = 32'h00000000;
    weight_b_mem[639] = 32'h00000000;
    weight_b_mem[640] = 32'h00000000;
    weight_b_mem[641] = 32'h00000000;
    weight_b_mem[642] = 32'h00000000;
    weight_b_mem[643] = 32'h00000000;
    weight_b_mem[644] = 32'h00000000;
    weight_b_mem[645] = 32'h00000000;
    weight_b_mem[646] = 32'h00000000;
    weight_b_mem[647] = 32'h00000000;
    weight_b_mem[648] = 32'h00000000;
    weight_b_mem[649] = 32'h00000000;
    weight_b_mem[650] = 32'h00000000;
    weight_b_mem[651] = 32'h00000000;
    weight_b_mem[652] = 32'h00000000;
    weight_b_mem[653] = 32'h00000000;
    weight_b_mem[654] = 32'h00000000;
    weight_b_mem[655] = 32'h00000000;
    weight_b_mem[656] = 32'h00000000;
    weight_b_mem[657] = 32'h00000000;
    weight_b_mem[658] = 32'h00000000;
    weight_b_mem[659] = 32'h00000000;
    weight_b_mem[660] = 32'h00000000;
    weight_b_mem[661] = 32'h00000000;
    weight_b_mem[662] = 32'h00000000;
    weight_b_mem[663] = 32'h00000000;
    weight_b_mem[664] = 32'h00000000;
    weight_b_mem[665] = 32'h00000000;
    weight_b_mem[666] = 32'h00000000;
    weight_b_mem[667] = 32'h00000000;
    weight_b_mem[668] = 32'h00000000;
    weight_b_mem[669] = 32'h00000000;
    weight_b_mem[670] = 32'h00000000;
    weight_b_mem[671] = 32'h00000000;
    weight_b_mem[672] = 32'h00000000;
    weight_b_mem[673] = 32'h00000000;
    weight_b_mem[674] = 32'h00000000;
    weight_b_mem[675] = 32'h00000000;
    weight_b_mem[676] = 32'h00000000;
    weight_b_mem[677] = 32'h00000000;
    weight_b_mem[678] = 32'h00000000;
    weight_b_mem[679] = 32'h00000000;
    weight_b_mem[680] = 32'h00000000;
    weight_b_mem[681] = 32'h00000000;
    weight_b_mem[682] = 32'h00000000;
    weight_b_mem[683] = 32'h00000000;
    weight_b_mem[684] = 32'h00000000;
    weight_b_mem[685] = 32'h00000000;
    weight_b_mem[686] = 32'h00000000;
    weight_b_mem[687] = 32'h00000000;
    weight_b_mem[688] = 32'h00000000;
    weight_b_mem[689] = 32'h00000000;
    weight_b_mem[690] = 32'h00000000;
    weight_b_mem[691] = 32'h00000000;
    weight_b_mem[692] = 32'h00000000;
    weight_b_mem[693] = 32'h00000000;
    weight_b_mem[694] = 32'h00000000;
    weight_b_mem[695] = 32'h00000000;
    weight_b_mem[696] = 32'h00000000;
    weight_b_mem[697] = 32'h00000000;
    weight_b_mem[698] = 32'h00000000;
    weight_b_mem[699] = 32'h00000000;
    weight_b_mem[700] = 32'h00000000;
    weight_b_mem[701] = 32'h00000000;
    weight_b_mem[702] = 32'h00000000;
    weight_b_mem[703] = 32'h00000000;
    weight_b_mem[704] = 32'h00000000;
    weight_b_mem[705] = 32'h00000000;
    weight_b_mem[706] = 32'h00000000;
    weight_b_mem[707] = 32'h00000000;
    weight_b_mem[708] = 32'h00000000;
    weight_b_mem[709] = 32'h00000000;
    weight_b_mem[710] = 32'h00000000;
    weight_b_mem[711] = 32'h00000000;
    weight_b_mem[712] = 32'h00000000;
    weight_b_mem[713] = 32'h00000000;
    weight_b_mem[714] = 32'h00000000;
    weight_b_mem[715] = 32'h00000000;
    weight_b_mem[716] = 32'h00000000;
    weight_b_mem[717] = 32'h00000000;
    weight_b_mem[718] = 32'h00000000;
    weight_b_mem[719] = 32'h00000000;
    weight_b_mem[720] = 32'h00000000;
    weight_b_mem[721] = 32'h00000000;
    weight_b_mem[722] = 32'h00000000;
    weight_b_mem[723] = 32'h00000000;
    weight_b_mem[724] = 32'h00000000;
    weight_b_mem[725] = 32'h00000000;
    weight_b_mem[726] = 32'h00000000;
    weight_b_mem[727] = 32'h00000000;
    weight_b_mem[728] = 32'h00000000;
    weight_b_mem[729] = 32'h00000000;
    weight_b_mem[730] = 32'h00000000;
    weight_b_mem[731] = 32'h00000000;
    weight_b_mem[732] = 32'h00000000;
    weight_b_mem[733] = 32'h00000000;
    weight_b_mem[734] = 32'h00000000;
    weight_b_mem[735] = 32'h00000000;
    weight_b_mem[736] = 32'h00000000;
    weight_b_mem[737] = 32'h00000000;
    weight_b_mem[738] = 32'h00000000;
    weight_b_mem[739] = 32'h00000000;
    weight_b_mem[740] = 32'h00000000;
    weight_b_mem[741] = 32'h00000000;
    weight_b_mem[742] = 32'h00000000;
    weight_b_mem[743] = 32'h00000000;
    weight_b_mem[744] = 32'h00000000;
    weight_b_mem[745] = 32'h00000000;
    weight_b_mem[746] = 32'h00000000;
    weight_b_mem[747] = 32'h00000000;
    weight_b_mem[748] = 32'h00000000;
    weight_b_mem[749] = 32'h00000000;
    weight_b_mem[750] = 32'h00000000;
    weight_b_mem[751] = 32'h00000000;
    weight_b_mem[752] = 32'h00000000;
    weight_b_mem[753] = 32'h00000000;
    weight_b_mem[754] = 32'h00000000;
    weight_b_mem[755] = 32'h00000000;
    weight_b_mem[756] = 32'h00000000;
    weight_b_mem[757] = 32'h00000000;
    weight_b_mem[758] = 32'h00000000;
    weight_b_mem[759] = 32'h00000000;
    weight_b_mem[760] = 32'h00000000;
    weight_b_mem[761] = 32'h00000000;
    weight_b_mem[762] = 32'h00000000;
    weight_b_mem[763] = 32'h00000000;
    weight_b_mem[764] = 32'h00000000;
    weight_b_mem[765] = 32'h00000000;
    weight_b_mem[766] = 32'h00000000;
    weight_b_mem[767] = 32'h00000000;
    weight_b_mem[768] = 32'h00000000;
    weight_b_mem[769] = 32'h00000000;
    weight_b_mem[770] = 32'h00000000;
    weight_b_mem[771] = 32'h00000000;
    weight_b_mem[772] = 32'h00000000;
    weight_b_mem[773] = 32'h00000000;
    weight_b_mem[774] = 32'h00000000;
    weight_b_mem[775] = 32'h00000000;
    weight_b_mem[776] = 32'h00000000;
    weight_b_mem[777] = 32'h00000000;
    weight_b_mem[778] = 32'h00000000;
    weight_b_mem[779] = 32'h00000000;
    weight_b_mem[780] = 32'h00000000;
    weight_b_mem[781] = 32'h00000000;
    weight_b_mem[782] = 32'h00000000;
    weight_b_mem[783] = 32'h00000000;
    weight_b_mem[784] = 32'h00000000;
    weight_b_mem[785] = 32'h00000000;
    weight_b_mem[786] = 32'h00000000;
    weight_b_mem[787] = 32'h00000000;
    weight_b_mem[788] = 32'h00000000;
    weight_b_mem[789] = 32'h00000000;
    weight_b_mem[790] = 32'h00000000;
    weight_b_mem[791] = 32'h00000000;
    weight_b_mem[792] = 32'h00000000;
    weight_b_mem[793] = 32'h00000000;
    weight_b_mem[794] = 32'h00000000;
    weight_b_mem[795] = 32'h00000000;
    weight_b_mem[796] = 32'h00000000;
    weight_b_mem[797] = 32'h00000000;
    weight_b_mem[798] = 32'h00000000;
    weight_b_mem[799] = 32'h00000000;
    weight_b_mem[800] = 32'h00000000;
    weight_b_mem[801] = 32'h00000000;
    weight_b_mem[802] = 32'h00000000;
    weight_b_mem[803] = 32'h00000000;
    weight_b_mem[804] = 32'h00000000;
    weight_b_mem[805] = 32'h00000000;
    weight_b_mem[806] = 32'h00000000;
    weight_b_mem[807] = 32'h00000000;
    weight_b_mem[808] = 32'h00000000;
    weight_b_mem[809] = 32'h00000000;
    weight_b_mem[810] = 32'h00000000;
    weight_b_mem[811] = 32'h00000000;
    weight_b_mem[812] = 32'h00000000;
    weight_b_mem[813] = 32'h00000000;
    weight_b_mem[814] = 32'h00000000;
    weight_b_mem[815] = 32'h00000000;
    weight_b_mem[816] = 32'h00000000;
    weight_b_mem[817] = 32'h00000000;
    weight_b_mem[818] = 32'h00000000;
    weight_b_mem[819] = 32'h00000000;
    weight_b_mem[820] = 32'h00000000;
    weight_b_mem[821] = 32'h00000000;
    weight_b_mem[822] = 32'h00000000;
    weight_b_mem[823] = 32'h00000000;
    weight_b_mem[824] = 32'h00000000;
    weight_b_mem[825] = 32'h00000000;
    weight_b_mem[826] = 32'h00000000;
    weight_b_mem[827] = 32'h00000000;
    weight_b_mem[828] = 32'h00000000;
    weight_b_mem[829] = 32'h00000000;
    weight_b_mem[830] = 32'h00000000;
    weight_b_mem[831] = 32'h00000000;
    weight_b_mem[832] = 32'h00000000;
    weight_b_mem[833] = 32'h00000000;
    weight_b_mem[834] = 32'h00000000;
    weight_b_mem[835] = 32'h00000000;
    weight_b_mem[836] = 32'h00000000;
    weight_b_mem[837] = 32'h00000000;
    weight_b_mem[838] = 32'h00000000;
    weight_b_mem[839] = 32'h00000000;
    weight_b_mem[840] = 32'h00000000;
    weight_b_mem[841] = 32'h00000000;
    weight_b_mem[842] = 32'h00000000;
    weight_b_mem[843] = 32'h00000000;
    weight_b_mem[844] = 32'h00000000;
    weight_b_mem[845] = 32'h00000000;
    weight_b_mem[846] = 32'h00000000;
    weight_b_mem[847] = 32'h00000000;
    weight_b_mem[848] = 32'h00000000;
    weight_b_mem[849] = 32'h00000000;
    weight_b_mem[850] = 32'h00000000;
    weight_b_mem[851] = 32'h00000000;
    weight_b_mem[852] = 32'h00000000;
    weight_b_mem[853] = 32'h00000000;
    weight_b_mem[854] = 32'h00000000;
    weight_b_mem[855] = 32'h00000000;
    weight_b_mem[856] = 32'h00000000;
    weight_b_mem[857] = 32'h00000000;
    weight_b_mem[858] = 32'h00000000;
    weight_b_mem[859] = 32'h00000000;
    weight_b_mem[860] = 32'h00000000;
    weight_b_mem[861] = 32'h00000000;
    weight_b_mem[862] = 32'h00000000;
    weight_b_mem[863] = 32'h00000000;
    weight_b_mem[864] = 32'h00000000;
    weight_b_mem[865] = 32'h00000000;
    weight_b_mem[866] = 32'h00000000;
    weight_b_mem[867] = 32'h00000000;
    weight_b_mem[868] = 32'h00000000;
    weight_b_mem[869] = 32'h00000000;
    weight_b_mem[870] = 32'h00000000;
    weight_b_mem[871] = 32'h00000000;
    weight_b_mem[872] = 32'h00000000;
    weight_b_mem[873] = 32'h00000000;
    weight_b_mem[874] = 32'h00000000;
    weight_b_mem[875] = 32'h00000000;
    weight_b_mem[876] = 32'h00000000;
    weight_b_mem[877] = 32'h00000000;
    weight_b_mem[878] = 32'h00000000;
    weight_b_mem[879] = 32'h00000000;
    weight_b_mem[880] = 32'h00000000;
    weight_b_mem[881] = 32'h00000000;
    weight_b_mem[882] = 32'h00000000;
    weight_b_mem[883] = 32'h00000000;
    weight_b_mem[884] = 32'h00000000;
    weight_b_mem[885] = 32'h00000000;
    weight_b_mem[886] = 32'h00000000;
    weight_b_mem[887] = 32'h00000000;
    weight_b_mem[888] = 32'h00000000;
    weight_b_mem[889] = 32'h00000000;
    weight_b_mem[890] = 32'h00000000;
    weight_b_mem[891] = 32'h00000000;
    weight_b_mem[892] = 32'h00000000;
    weight_b_mem[893] = 32'h00000000;
    weight_b_mem[894] = 32'h00000000;
    weight_b_mem[895] = 32'h00000000;
    weight_b_mem[896] = 32'h00000000;
    weight_b_mem[897] = 32'h00000000;
    weight_b_mem[898] = 32'h00000000;
    weight_b_mem[899] = 32'h00000000;
    weight_b_mem[900] = 32'h00000000;
    weight_b_mem[901] = 32'h00000000;
    weight_b_mem[902] = 32'h00000000;
    weight_b_mem[903] = 32'h00000000;
    weight_b_mem[904] = 32'h00000000;
    weight_b_mem[905] = 32'h00000000;
    weight_b_mem[906] = 32'h00000000;
    weight_b_mem[907] = 32'h00000000;
    weight_b_mem[908] = 32'h00000000;
    weight_b_mem[909] = 32'h00000000;
    weight_b_mem[910] = 32'h00000000;
    weight_b_mem[911] = 32'h00000000;
    weight_b_mem[912] = 32'h00000000;
    weight_b_mem[913] = 32'h00000000;
    weight_b_mem[914] = 32'h00000000;
    weight_b_mem[915] = 32'h00000000;
    weight_b_mem[916] = 32'h00000000;
    weight_b_mem[917] = 32'h00000000;
    weight_b_mem[918] = 32'h00000000;
    weight_b_mem[919] = 32'h00000000;
    weight_b_mem[920] = 32'h00000000;
    weight_b_mem[921] = 32'h00000000;
    weight_b_mem[922] = 32'h00000000;
    weight_b_mem[923] = 32'h00000000;
    weight_b_mem[924] = 32'h00000000;
    weight_b_mem[925] = 32'h00000000;
    weight_b_mem[926] = 32'h00000000;
    weight_b_mem[927] = 32'h00000000;
    weight_b_mem[928] = 32'h00000000;
    weight_b_mem[929] = 32'h00000000;
    weight_b_mem[930] = 32'h00000000;
    weight_b_mem[931] = 32'h00000000;
    weight_b_mem[932] = 32'h00000000;
    weight_b_mem[933] = 32'h00000000;
    weight_b_mem[934] = 32'h00000000;
    weight_b_mem[935] = 32'h00000000;
    weight_b_mem[936] = 32'h00000000;
    weight_b_mem[937] = 32'h00000000;
    weight_b_mem[938] = 32'h00000000;
    weight_b_mem[939] = 32'h00000000;
    weight_b_mem[940] = 32'h00000000;
    weight_b_mem[941] = 32'h00000000;
    weight_b_mem[942] = 32'h00000000;
    weight_b_mem[943] = 32'h00000000;
    weight_b_mem[944] = 32'h00000000;
    weight_b_mem[945] = 32'h00000000;
    weight_b_mem[946] = 32'h00000000;
    weight_b_mem[947] = 32'h00000000;
    weight_b_mem[948] = 32'h00000000;
    weight_b_mem[949] = 32'h00000000;
    weight_b_mem[950] = 32'h00000000;
    weight_b_mem[951] = 32'h00000000;
    weight_b_mem[952] = 32'h00000000;
    weight_b_mem[953] = 32'h00000000;
    weight_b_mem[954] = 32'h00000000;
    weight_b_mem[955] = 32'h00000000;
    weight_b_mem[956] = 32'h00000000;
    weight_b_mem[957] = 32'h00000000;
    weight_b_mem[958] = 32'h00000000;
    weight_b_mem[959] = 32'h00000000;
    weight_b_mem[960] = 32'h00000000;
    weight_b_mem[961] = 32'h00000000;
    weight_b_mem[962] = 32'h00000000;
    weight_b_mem[963] = 32'h00000000;
    weight_b_mem[964] = 32'h00000000;
    weight_b_mem[965] = 32'h00000000;
    weight_b_mem[966] = 32'h00000000;
    weight_b_mem[967] = 32'h00000000;
    weight_b_mem[968] = 32'h00000000;
    weight_b_mem[969] = 32'h00000000;
    weight_b_mem[970] = 32'h00000000;
    weight_b_mem[971] = 32'h00000000;
    weight_b_mem[972] = 32'h00000000;
    weight_b_mem[973] = 32'h00000000;
    weight_b_mem[974] = 32'h00000000;
    weight_b_mem[975] = 32'h00000000;
    weight_b_mem[976] = 32'h00000000;
    weight_b_mem[977] = 32'h00000000;
    weight_b_mem[978] = 32'h00000000;
    weight_b_mem[979] = 32'h00000000;
    weight_b_mem[980] = 32'h00000000;
    weight_b_mem[981] = 32'h00000000;
    weight_b_mem[982] = 32'h00000000;
    weight_b_mem[983] = 32'h00000000;
    weight_b_mem[984] = 32'h00000000;
    weight_b_mem[985] = 32'h00000000;
    weight_b_mem[986] = 32'h00000000;
    weight_b_mem[987] = 32'h00000000;
    weight_b_mem[988] = 32'h00000000;
    weight_b_mem[989] = 32'h00000000;
    weight_b_mem[990] = 32'h00000000;
    weight_b_mem[991] = 32'h00000000;
    weight_b_mem[992] = 32'h00000000;
    weight_b_mem[993] = 32'h00000000;
    weight_b_mem[994] = 32'h00000000;
    weight_b_mem[995] = 32'h00000000;
    weight_b_mem[996] = 32'h00000000;
    weight_b_mem[997] = 32'h00000000;
    weight_b_mem[998] = 32'h00000000;
    weight_b_mem[999] = 32'h00000000;
    weight_b_mem[1000] = 32'h00000000;
    weight_b_mem[1001] = 32'h00000000;
    weight_b_mem[1002] = 32'h00000000;
    weight_b_mem[1003] = 32'h00000000;
    weight_b_mem[1004] = 32'h00000000;
    weight_b_mem[1005] = 32'h00000000;
    weight_b_mem[1006] = 32'h00000000;
    weight_b_mem[1007] = 32'h00000000;
    weight_b_mem[1008] = 32'h00000000;
    weight_b_mem[1009] = 32'h00000000;
    weight_b_mem[1010] = 32'h00000000;
    weight_b_mem[1011] = 32'h00000000;
    weight_b_mem[1012] = 32'h00000000;
    weight_b_mem[1013] = 32'h00000000;
    weight_b_mem[1014] = 32'h00000000;
    weight_b_mem[1015] = 32'h00000000;
    weight_b_mem[1016] = 32'h00000000;
    weight_b_mem[1017] = 32'h00000000;
    weight_b_mem[1018] = 32'h00000000;
    weight_b_mem[1019] = 32'h00000000;
    weight_b_mem[1020] = 32'h00000000;
    weight_b_mem[1021] = 32'h00000000;
    weight_b_mem[1022] = 32'h00000000;
    weight_b_mem[1023] = 32'h00000000;
    weight_b_mem[1024] = 32'h00000000;
    weight_b_mem[1025] = 32'h00000000;
    weight_b_mem[1026] = 32'h00000000;
    weight_b_mem[1027] = 32'h00000000;
    weight_b_mem[1028] = 32'h00000000;
    weight_b_mem[1029] = 32'h00000000;
    weight_b_mem[1030] = 32'h00000000;
    weight_b_mem[1031] = 32'h00000000;
    weight_b_mem[1032] = 32'h00000000;
    weight_b_mem[1033] = 32'h00000000;
    weight_b_mem[1034] = 32'h00000000;
    weight_b_mem[1035] = 32'h00000000;
    weight_b_mem[1036] = 32'h00000000;
    weight_b_mem[1037] = 32'h00000000;
    weight_b_mem[1038] = 32'h00000000;
    weight_b_mem[1039] = 32'h00000000;
    weight_b_mem[1040] = 32'h00000000;
    weight_b_mem[1041] = 32'h00000000;
    weight_b_mem[1042] = 32'h00000000;
    weight_b_mem[1043] = 32'h00000000;
    weight_b_mem[1044] = 32'h00000000;
    weight_b_mem[1045] = 32'h00000000;
    weight_b_mem[1046] = 32'h00000000;
    weight_b_mem[1047] = 32'h00000000;
    weight_b_mem[1048] = 32'h00000000;
    weight_b_mem[1049] = 32'h00000000;
    weight_b_mem[1050] = 32'h00000000;
    weight_b_mem[1051] = 32'h00000000;
    weight_b_mem[1052] = 32'h00000000;
    weight_b_mem[1053] = 32'h00000000;
    weight_b_mem[1054] = 32'h00000000;
    weight_b_mem[1055] = 32'h00000000;
    weight_b_mem[1056] = 32'h00000000;
    weight_b_mem[1057] = 32'h00000000;
    weight_b_mem[1058] = 32'h00000000;
    weight_b_mem[1059] = 32'h00000000;
    weight_b_mem[1060] = 32'h00000000;
    weight_b_mem[1061] = 32'h00000000;
    weight_b_mem[1062] = 32'h00000000;
    weight_b_mem[1063] = 32'h00000000;
    weight_b_mem[1064] = 32'h00000000;
    weight_b_mem[1065] = 32'h00000000;
    weight_b_mem[1066] = 32'h00000000;
    weight_b_mem[1067] = 32'h00000000;
    weight_b_mem[1068] = 32'h00000000;
    weight_b_mem[1069] = 32'h00000000;
    weight_b_mem[1070] = 32'h00000000;
    weight_b_mem[1071] = 32'h00000000;
    weight_b_mem[1072] = 32'h00000000;
    weight_b_mem[1073] = 32'h00000000;
    weight_b_mem[1074] = 32'h00000000;
    weight_b_mem[1075] = 32'h00000000;
    weight_b_mem[1076] = 32'h00000000;
    weight_b_mem[1077] = 32'h00000000;
    weight_b_mem[1078] = 32'h00000000;
    weight_b_mem[1079] = 32'h00000000;
    weight_b_mem[1080] = 32'h00000000;
    weight_b_mem[1081] = 32'h00000000;
    weight_b_mem[1082] = 32'h00000000;
    weight_b_mem[1083] = 32'h00000000;
    weight_b_mem[1084] = 32'h00000000;
    weight_b_mem[1085] = 32'h00000000;
    weight_b_mem[1086] = 32'h00000000;
    weight_b_mem[1087] = 32'h00000000;
    weight_b_mem[1088] = 32'h00000000;
    weight_b_mem[1089] = 32'h00000000;
    weight_b_mem[1090] = 32'h00000000;
    weight_b_mem[1091] = 32'h00000000;
    weight_b_mem[1092] = 32'h00000000;
    weight_b_mem[1093] = 32'h00000000;
    weight_b_mem[1094] = 32'h00000000;
    weight_b_mem[1095] = 32'h00000000;
    weight_b_mem[1096] = 32'h00000000;
    weight_b_mem[1097] = 32'h00000000;
    weight_b_mem[1098] = 32'h00000000;
    weight_b_mem[1099] = 32'h00000000;
    weight_b_mem[1100] = 32'h00000000;
    weight_b_mem[1101] = 32'h00000000;
    weight_b_mem[1102] = 32'h00000000;
    weight_b_mem[1103] = 32'h00000000;
    weight_b_mem[1104] = 32'h00000000;
    weight_b_mem[1105] = 32'h00000000;
    weight_b_mem[1106] = 32'h00000000;
    weight_b_mem[1107] = 32'h00000000;
    weight_b_mem[1108] = 32'h00000000;
    weight_b_mem[1109] = 32'h00000000;
    weight_b_mem[1110] = 32'h00000000;
    weight_b_mem[1111] = 32'h00000000;
    weight_b_mem[1112] = 32'h00000000;
    weight_b_mem[1113] = 32'h00000000;
    weight_b_mem[1114] = 32'h00000000;
    weight_b_mem[1115] = 32'h00000000;
    weight_b_mem[1116] = 32'h00000000;
    weight_b_mem[1117] = 32'h00000000;
    weight_b_mem[1118] = 32'h00000000;
    weight_b_mem[1119] = 32'h00000000;
    weight_b_mem[1120] = 32'h00000000;
    weight_b_mem[1121] = 32'h00000000;
    weight_b_mem[1122] = 32'h00000000;
    weight_b_mem[1123] = 32'h00000000;
    weight_b_mem[1124] = 32'h00000000;
    weight_b_mem[1125] = 32'h00000000;
    weight_b_mem[1126] = 32'h00000000;
    weight_b_mem[1127] = 32'h00000000;
    weight_b_mem[1128] = 32'h00000000;
    weight_b_mem[1129] = 32'h00000000;
    weight_b_mem[1130] = 32'h00000000;
    weight_b_mem[1131] = 32'h00000000;
    weight_b_mem[1132] = 32'h00000000;
    weight_b_mem[1133] = 32'h00000000;
    weight_b_mem[1134] = 32'h00000000;
    weight_b_mem[1135] = 32'h00000000;
    weight_b_mem[1136] = 32'h00000000;
    weight_b_mem[1137] = 32'h00000000;
    weight_b_mem[1138] = 32'h00000000;
    weight_b_mem[1139] = 32'h00000000;
    weight_b_mem[1140] = 32'h00000000;
    weight_b_mem[1141] = 32'h00000000;
    weight_b_mem[1142] = 32'h00000000;
    weight_b_mem[1143] = 32'h00000000;
    weight_b_mem[1144] = 32'h00000000;
    weight_b_mem[1145] = 32'h00000000;
    weight_b_mem[1146] = 32'h00000000;
    weight_b_mem[1147] = 32'h00000000;
    weight_b_mem[1148] = 32'h00000000;
    weight_b_mem[1149] = 32'h00000000;
    weight_b_mem[1150] = 32'h00000000;
    weight_b_mem[1151] = 32'h00000000;
    weight_b_mem[1152] = 32'h00000000;
    weight_b_mem[1153] = 32'h00000000;
    weight_b_mem[1154] = 32'h00000000;
    weight_b_mem[1155] = 32'h00000000;
    weight_b_mem[1156] = 32'h00000000;
    weight_b_mem[1157] = 32'h00000000;
    weight_b_mem[1158] = 32'h00000000;
    weight_b_mem[1159] = 32'h00000000;
    weight_b_mem[1160] = 32'h00000000;
    weight_b_mem[1161] = 32'h00000000;
    weight_b_mem[1162] = 32'h00000000;
    weight_b_mem[1163] = 32'h00000000;
    weight_b_mem[1164] = 32'h00000000;
    weight_b_mem[1165] = 32'h00000000;
    weight_b_mem[1166] = 32'h00000000;
    weight_b_mem[1167] = 32'h00000000;
    weight_b_mem[1168] = 32'h00000000;
    weight_b_mem[1169] = 32'h00000000;
    weight_b_mem[1170] = 32'h00000000;
    weight_b_mem[1171] = 32'h00000000;
    weight_b_mem[1172] = 32'h00000000;
    weight_b_mem[1173] = 32'h00000000;
    weight_b_mem[1174] = 32'h00000000;
    weight_b_mem[1175] = 32'h00000000;
    weight_b_mem[1176] = 32'h00000000;
    weight_b_mem[1177] = 32'h00000000;
    weight_b_mem[1178] = 32'h00000000;
    weight_b_mem[1179] = 32'h00000000;
    weight_b_mem[1180] = 32'h00000000;
    weight_b_mem[1181] = 32'h00000000;
    weight_b_mem[1182] = 32'h00000000;
    weight_b_mem[1183] = 32'h00000000;
    weight_b_mem[1184] = 32'h00000000;
    weight_b_mem[1185] = 32'h00000000;
    weight_b_mem[1186] = 32'h00000000;
    weight_b_mem[1187] = 32'h00000000;
    weight_b_mem[1188] = 32'h00000000;
    weight_b_mem[1189] = 32'h00000000;
    weight_b_mem[1190] = 32'h00000000;
    weight_b_mem[1191] = 32'h00000000;
    weight_b_mem[1192] = 32'h00000000;
    weight_b_mem[1193] = 32'h00000000;
    weight_b_mem[1194] = 32'h00000000;
    weight_b_mem[1195] = 32'h00000000;
    weight_b_mem[1196] = 32'h00000000;
    weight_b_mem[1197] = 32'h00000000;
    weight_b_mem[1198] = 32'h00000000;
    weight_b_mem[1199] = 32'h00000000;
    weight_b_mem[1200] = 32'h00000000;
    weight_b_mem[1201] = 32'h00000000;
    weight_b_mem[1202] = 32'h00000000;
    weight_b_mem[1203] = 32'h00000000;
    weight_b_mem[1204] = 32'h00000000;
    weight_b_mem[1205] = 32'h00000000;
    weight_b_mem[1206] = 32'h00000000;
    weight_b_mem[1207] = 32'h00000000;
    weight_b_mem[1208] = 32'h00000000;
    weight_b_mem[1209] = 32'h00000000;
    weight_b_mem[1210] = 32'h00000000;
    weight_b_mem[1211] = 32'h00000000;
    weight_b_mem[1212] = 32'h00000000;
    weight_b_mem[1213] = 32'h00000000;
    weight_b_mem[1214] = 32'h00000000;
    weight_b_mem[1215] = 32'h00000000;
    weight_b_mem[1216] = 32'h00000000;
    weight_b_mem[1217] = 32'h00000000;
    weight_b_mem[1218] = 32'h00000000;
    weight_b_mem[1219] = 32'h00000000;
    weight_b_mem[1220] = 32'h00000000;
    weight_b_mem[1221] = 32'h00000000;
    weight_b_mem[1222] = 32'h00000000;
    weight_b_mem[1223] = 32'h00000000;
    weight_b_mem[1224] = 32'h00000000;
    weight_b_mem[1225] = 32'h00000000;
    weight_b_mem[1226] = 32'h00000000;
    weight_b_mem[1227] = 32'h00000000;
    weight_b_mem[1228] = 32'h00000000;
    weight_b_mem[1229] = 32'h00000000;
    weight_b_mem[1230] = 32'h00000000;
    weight_b_mem[1231] = 32'h00000000;
    weight_b_mem[1232] = 32'h00000000;
    weight_b_mem[1233] = 32'h00000000;
    weight_b_mem[1234] = 32'h00000000;
    weight_b_mem[1235] = 32'h00000000;
    weight_b_mem[1236] = 32'h00000000;
    weight_b_mem[1237] = 32'h00000000;
    weight_b_mem[1238] = 32'h00000000;
    weight_b_mem[1239] = 32'h00000000;
    weight_b_mem[1240] = 32'h00000000;
    weight_b_mem[1241] = 32'h00000000;
    weight_b_mem[1242] = 32'h00000000;
    weight_b_mem[1243] = 32'h00000000;
    weight_b_mem[1244] = 32'h00000000;
    weight_b_mem[1245] = 32'h00000000;
    weight_b_mem[1246] = 32'h00000000;
    weight_b_mem[1247] = 32'h00000000;
    weight_b_mem[1248] = 32'h00000000;
    weight_b_mem[1249] = 32'h00000000;
    weight_b_mem[1250] = 32'h00000000;
    weight_b_mem[1251] = 32'h00000000;
    weight_b_mem[1252] = 32'h00000000;
    weight_b_mem[1253] = 32'h00000000;
    weight_b_mem[1254] = 32'h00000000;
    weight_b_mem[1255] = 32'h00000000;
    weight_b_mem[1256] = 32'h00000000;
    weight_b_mem[1257] = 32'h00000000;
    weight_b_mem[1258] = 32'h00000000;
    weight_b_mem[1259] = 32'h00000000;
    weight_b_mem[1260] = 32'h00000000;
    weight_b_mem[1261] = 32'h00000000;
    weight_b_mem[1262] = 32'h00000000;
    weight_b_mem[1263] = 32'h00000000;
    weight_b_mem[1264] = 32'h00000000;
    weight_b_mem[1265] = 32'h00000000;
    weight_b_mem[1266] = 32'h00000000;
    weight_b_mem[1267] = 32'h00000000;
    weight_b_mem[1268] = 32'h00000000;
    weight_b_mem[1269] = 32'h00000000;
    weight_b_mem[1270] = 32'h00000000;
    weight_b_mem[1271] = 32'h00000000;
    weight_b_mem[1272] = 32'h00000000;
    weight_b_mem[1273] = 32'h00000000;
    weight_b_mem[1274] = 32'h00000000;
    weight_b_mem[1275] = 32'h00000000;
    weight_b_mem[1276] = 32'h00000000;
    weight_b_mem[1277] = 32'h00000000;
    weight_b_mem[1278] = 32'h00000000;
    weight_b_mem[1279] = 32'h00000000;
    weight_b_mem[1280] = 32'h00000000;
    weight_b_mem[1281] = 32'h00000000;
    weight_b_mem[1282] = 32'h00000000;
end
