// sine_lut.v — Quarter-wave sine lookup table for SIREN activation
//
// Computes sin(angle) for Q4.28 fixed-point inputs and outputs.
// Uses 256-entry quarter-wave table with quadrant reconstruction.
//
// Input:  angle in Q4.28 radians (any value, reduced mod 2*pi)
// Output: sin(angle) in Q4.28 (range [-1, +1])
//
// Latency: 2 cycles (registered input + registered output)
//
// For SIREN networks, the activation is sin(omega * x) where omega
// is typically 30.0 for the first layer and 1.0 for hidden layers.
// The omega scaling is done in the MLP core before calling this LUT.

`timescale 1ns / 1ps

module sine_lut #(
    parameter WIDTH = 32,
    parameter FRAC  = 28
)(
    input  wire                    clk,
    input  wire signed [WIDTH-1:0] angle,   // Q4.28 radians
    output reg  signed [WIDTH-1:0] result   // Q4.28 sin(angle)
);

    // =========================================================
    // Constants in Q4.28
    // =========================================================
    // pi   = 3.14159265... * 2^28 = 843314857  = 32'h3243_F6A9
    // 2*pi = 6.28318530... * 2^28 = 1686629713 = 32'h6487_ED51
    // pi/2 = 1.57079632... * 2^28 = 421657428  = 32'h1921_FB54
    localparam signed [WIDTH-1:0] TWO_PI  = 32'sh6487_ED51;
    localparam signed [WIDTH-1:0] PI      = 32'sh3243_F6A9;
    localparam signed [WIDTH-1:0] HALF_PI = 32'sh1921_FB54;

    // =========================================================
    // Quarter-wave sine table: 256 entries for [0, pi/2)
    // =========================================================
    // Entry k = sin(k * pi/2 / 256) in Q4.28
    // sin(0) = 0, sin(pi/2) = 1.0 = 0x10000000
    //
    // Generated by: round(sin(k * pi / 512) * 2^28) for k=0..255
    reg signed [WIDTH-1:0] sine_table [0:255];

    initial begin
        sine_table[  0] = 32'sh00000000; sine_table[  1] = 32'sh00C90F88;
        sine_table[  2] = 32'sh01921D20; sine_table[  3] = 32'sh025B26D7;
        sine_table[  4] = 32'sh03242ABF; sine_table[  5] = 32'sh03ED26E6;
        sine_table[  6] = 32'sh04B6195D; sine_table[  7] = 32'sh057F0035;
        sine_table[  8] = 32'sh0647D97C; sine_table[  9] = 32'sh0710A345;
        sine_table[ 10] = 32'sh07D95B9E; sine_table[ 11] = 32'sh08A2009A;
        sine_table[ 12] = 32'sh096A9049; sine_table[ 13] = 32'sh0A3308BD;
        sine_table[ 14] = 32'sh0AFB6805; sine_table[ 15] = 32'sh0BC3AC35;
        sine_table[ 16] = 32'sh0C8BD35E; sine_table[ 17] = 32'sh0D53DB92;
        sine_table[ 18] = 32'sh0E1BC2E4; sine_table[ 19] = 32'sh0EE38766;
        sine_table[ 20] = 32'sh0FAB272B; sine_table[ 21] = 32'sh1072A048;
        sine_table[ 22] = 32'sh1139F0CF; sine_table[ 23] = 32'sh120116D5;
        sine_table[ 24] = 32'sh12C8106F; sine_table[ 25] = 32'sh138EDBB1;
        sine_table[ 26] = 32'sh145576B1; sine_table[ 27] = 32'sh151BDF86;
        sine_table[ 28] = 32'sh15E21445; sine_table[ 29] = 32'sh16A81305;
        sine_table[ 30] = 32'sh176DD9DE; sine_table[ 31] = 32'sh183366E9;
        sine_table[ 32] = 32'sh18F8B83C; sine_table[ 33] = 32'sh19BDCBF3;
        sine_table[ 34] = 32'sh1A82A026; sine_table[ 35] = 32'sh1B4732EF;
        sine_table[ 36] = 32'sh1C0B826A; sine_table[ 37] = 32'sh1CCF8CB3;
        sine_table[ 38] = 32'sh1D934FE5; sine_table[ 39] = 32'sh1E56CA1E;
        sine_table[ 40] = 32'sh1F19F97B; sine_table[ 41] = 32'sh1FDCDC1B;
        sine_table[ 42] = 32'sh209F701C; sine_table[ 43] = 32'sh2161B3A0;
        sine_table[ 44] = 32'sh2223A4C5; sine_table[ 45] = 32'sh22E541AF;
        sine_table[ 46] = 32'sh23A6887F; sine_table[ 47] = 32'sh24677758;
        sine_table[ 48] = 32'sh25280C5E; sine_table[ 49] = 32'sh25E845B6;
        sine_table[ 50] = 32'sh26A82186; sine_table[ 51] = 32'sh27679DF4;
        sine_table[ 52] = 32'sh2826B928; sine_table[ 53] = 32'sh28E5714B;
        sine_table[ 54] = 32'sh29A3C485; sine_table[ 55] = 32'sh2A61B101;
        sine_table[ 56] = 32'sh2B1F34EB; sine_table[ 57] = 32'sh2BDC4E6F;
        sine_table[ 58] = 32'sh2C98FBBA; sine_table[ 59] = 32'sh2D553AFB;
        sine_table[ 60] = 32'sh2E110A62; sine_table[ 61] = 32'sh2ECC681E;
        sine_table[ 62] = 32'sh2F875262; sine_table[ 63] = 32'sh3041C761;
        sine_table[ 64] = 32'sh30FBC54D; sine_table[ 65] = 32'sh31B54A5E;
        sine_table[ 66] = 32'sh326E54C7; sine_table[ 67] = 32'sh3326E2C3;
        sine_table[ 68] = 32'sh33DEF287; sine_table[ 69] = 32'sh3496824F;
        sine_table[ 70] = 32'sh354D9057; sine_table[ 71] = 32'sh36041AD9;
        sine_table[ 72] = 32'sh36BA2014; sine_table[ 73] = 32'sh376F9E46;
        sine_table[ 74] = 32'sh382493B0; sine_table[ 75] = 32'sh38D8FE93;
        sine_table[ 76] = 32'sh398CDD32; sine_table[ 77] = 32'sh3A402DD2;
        sine_table[ 78] = 32'sh3AF2EEB7; sine_table[ 79] = 32'sh3BA51E29;
        sine_table[ 80] = 32'sh3C56BA70; sine_table[ 81] = 32'sh3D07C1D6;
        sine_table[ 82] = 32'sh3DB832A6; sine_table[ 83] = 32'sh3E680B2C;
        sine_table[ 84] = 32'sh3F1749B8; sine_table[ 85] = 32'sh3FC5EC98;
        sine_table[ 86] = 32'sh4073F21D; sine_table[ 87] = 32'sh4121589B;
        sine_table[ 88] = 32'sh41CE1E65; sine_table[ 89] = 32'sh427A41D0;
        sine_table[ 90] = 32'sh4325C135; sine_table[ 91] = 32'sh43D09AED;
        sine_table[ 92] = 32'sh447ACD50; sine_table[ 93] = 32'sh452456BD;
        sine_table[ 94] = 32'sh45CD358F; sine_table[ 95] = 32'sh46756828;
        sine_table[ 96] = 32'sh471CECE7; sine_table[ 97] = 32'sh47C3C22F;
        sine_table[ 98] = 32'sh4869E665; sine_table[ 99] = 32'sh490F57EE;
        sine_table[100] = 32'sh49B41533; sine_table[101] = 32'sh4A581C9E;
        sine_table[102] = 32'sh4AFB6C98; sine_table[103] = 32'sh4B9E0390;
        sine_table[104] = 32'sh4C3FDFF4; sine_table[105] = 32'sh4CE10034;
        sine_table[106] = 32'sh4D8162C4; sine_table[107] = 32'sh4E210617;
        sine_table[108] = 32'sh4EBFE8A5; sine_table[109] = 32'sh4F5E08E3;
        sine_table[110] = 32'sh4FFB654D; sine_table[111] = 32'sh5097FC5E;
        sine_table[112] = 32'sh5133CC94; sine_table[113] = 32'sh51CED46E;
        sine_table[114] = 32'sh5269126E; sine_table[115] = 32'sh53028518;
        sine_table[116] = 32'sh539B2AF0; sine_table[117] = 32'sh5433027D;
        sine_table[118] = 32'sh54CA0A4B; sine_table[119] = 32'sh556040E2;
        sine_table[120] = 32'sh55F5A4D2; sine_table[121] = 32'sh568A34A9;
        sine_table[122] = 32'sh571DEEFA; sine_table[123] = 32'sh57B0D256;
        sine_table[124] = 32'sh5842DD54; sine_table[125] = 32'sh58D40E8C;
        sine_table[126] = 32'sh59646498; sine_table[127] = 32'sh59F3DE12;
        sine_table[128] = 32'sh5A82799A; sine_table[129] = 32'sh5B1035CF;
        sine_table[130] = 32'sh5B9D1154; sine_table[131] = 32'sh5C290ACC;
        sine_table[132] = 32'sh5CB420E0; sine_table[133] = 32'sh5D3E5237;
        sine_table[134] = 32'sh5DC79D7C; sine_table[135] = 32'sh5E50015D;
        sine_table[136] = 32'sh5ED77C8A; sine_table[137] = 32'sh5F5E0DB3;
        sine_table[138] = 32'sh5FE3B38D; sine_table[139] = 32'sh60686CCF;
        sine_table[140] = 32'sh60EC3830; sine_table[141] = 32'sh616F146C;
        sine_table[142] = 32'sh61F1003F; sine_table[143] = 32'sh6271FA69;
        sine_table[144] = 32'sh62F201AC; sine_table[145] = 32'sh637114CC;
        sine_table[146] = 32'sh63EF3290; sine_table[147] = 32'sh646C59BF;
        sine_table[148] = 32'sh64E88926; sine_table[149] = 32'sh6563BF92;
        sine_table[150] = 32'sh65DDFBD3; sine_table[151] = 32'sh66573CBB;
        sine_table[152] = 32'sh66CF8120; sine_table[153] = 32'sh6746C7D8;
        sine_table[154] = 32'sh67BD0FBD; sine_table[155] = 32'sh683257AB;
        sine_table[156] = 32'sh68A69E81; sine_table[157] = 32'sh6919E320;
        sine_table[158] = 32'sh698C246C; sine_table[159] = 32'sh69FD614A;
        sine_table[160] = 32'sh6A6D98A4; sine_table[161] = 32'sh6ADCC964;
        sine_table[162] = 32'sh6B4AF279; sine_table[163] = 32'sh6BB812D1;
        sine_table[164] = 32'sh6C242960; sine_table[165] = 32'sh6C8F351C;
        sine_table[166] = 32'sh6CF934FC; sine_table[167] = 32'sh6D6227FA;
        sine_table[168] = 32'sh6DCA0D14; sine_table[169] = 32'sh6E30E34A;
        sine_table[170] = 32'sh6E96A99D; sine_table[171] = 32'sh6EFB5F12;
        sine_table[172] = 32'sh6F5F02B2; sine_table[173] = 32'sh6FC19385;
        sine_table[174] = 32'sh70231099; sine_table[175] = 32'sh708378FF;
        sine_table[176] = 32'sh70E2CBC6; sine_table[177] = 32'sh71410805;
        sine_table[178] = 32'sh719E2CD2; sine_table[179] = 32'sh71FA3949;
        sine_table[180] = 32'sh72552C85; sine_table[181] = 32'sh72AF05A7;
        sine_table[182] = 32'sh7307C3D0; sine_table[183] = 32'sh735F6626;
        sine_table[184] = 32'sh73B5EBD1; sine_table[185] = 32'sh740B53FB;
        sine_table[186] = 32'sh745F9DD1; sine_table[187] = 32'sh74B2C884;
        sine_table[188] = 32'sh7504D345; sine_table[189] = 32'sh7555BD4C;
        sine_table[190] = 32'sh75A585CF; sine_table[191] = 32'sh75F42C0B;
        sine_table[192] = 32'sh7641AF3D; sine_table[193] = 32'sh768E0EA6;
        sine_table[194] = 32'sh76D94989; sine_table[195] = 32'sh77235F2D;
        sine_table[196] = 32'sh776C4EDB; sine_table[197] = 32'sh77B417DF;
        sine_table[198] = 32'sh77FAB989; sine_table[199] = 32'sh78403329;
        sine_table[200] = 32'sh78848414; sine_table[201] = 32'sh78C7ABA2;
        sine_table[202] = 32'sh7909A92D; sine_table[203] = 32'sh794A7C12;
        sine_table[204] = 32'sh798A23B1; sine_table[205] = 32'sh79C89F6E;
        sine_table[206] = 32'sh7A05EEAD; sine_table[207] = 32'sh7A4210D8;
        sine_table[208] = 32'sh7A7D055B; sine_table[209] = 32'sh7AB6CBA4;
        sine_table[210] = 32'sh7AEF6323; sine_table[211] = 32'sh7B26CB4F;
        sine_table[212] = 32'sh7B5D039E; sine_table[213] = 32'sh7B920B89;
        sine_table[214] = 32'sh7BC5E290; sine_table[215] = 32'sh7BF88830;
        sine_table[216] = 32'sh7C29FBEE; sine_table[217] = 32'sh7C5A3D50;
        sine_table[218] = 32'sh7C894BDE; sine_table[219] = 32'sh7CB72724;
        sine_table[220] = 32'sh7CE3CEB2; sine_table[221] = 32'sh7D0F4218;
        sine_table[222] = 32'sh7D3980EC; sine_table[223] = 32'sh7D628AC6;
        sine_table[224] = 32'sh7D8A5F40; sine_table[225] = 32'sh7DB0FDF8;
        sine_table[226] = 32'sh7DD6668F; sine_table[227] = 32'sh7DFA98A8;
        sine_table[228] = 32'sh7E1D93EA; sine_table[229] = 32'sh7E3F57FF;
        sine_table[230] = 32'sh7E5FE493; sine_table[231] = 32'sh7E7F3957;
        sine_table[232] = 32'sh7E9D55FC; sine_table[233] = 32'sh7EBA3A39;
        sine_table[234] = 32'sh7ED5E5C6; sine_table[235] = 32'sh7EF05860;
        sine_table[236] = 32'sh7F0991C4; sine_table[237] = 32'sh7F2191B4;
        sine_table[238] = 32'sh7F3857F6; sine_table[239] = 32'sh7F4DE451;
        sine_table[240] = 32'sh7F62368F; sine_table[241] = 32'sh7F754E80;
        sine_table[242] = 32'sh7F872BF3; sine_table[243] = 32'sh7F97CEBD;
        sine_table[244] = 32'sh7FA736B4; sine_table[245] = 32'sh7FB563B3;
        sine_table[246] = 32'sh7FC25596; sine_table[247] = 32'sh7FCE0C3E;
        sine_table[248] = 32'sh7FD8878E; sine_table[249] = 32'sh7FE1C76B;
        sine_table[250] = 32'sh7FE9CBC0; sine_table[251] = 32'sh7FF09478;
        sine_table[252] = 32'sh7FF62182; sine_table[253] = 32'sh7FFA72D1;
        sine_table[254] = 32'sh7FFD885A; sine_table[255] = 32'sh7FFF6217;
    end

    // =========================================================
    // Stage 1: Reduce angle mod 2*pi, determine quadrant
    // =========================================================
    // We need angle in [0, 2*pi). For the quarter-wave approach:
    //   quadrant 0: [0, pi/2)      → table[idx]
    //   quadrant 1: [pi/2, pi)     → table[255-idx]
    //   quadrant 2: [pi, 3pi/2)    → -table[idx]
    //   quadrant 3: [3pi/2, 2pi)   → -table[255-idx]

    // Modular reduction: we use the fractional bits after dividing by 2*pi.
    // angle / (2*pi) gives us the fractional position in the cycle.
    // We approximate by using the upper bits of (angle * (1/(2*pi))).
    //
    // Simpler approach: since we only need 256 entries per quadrant,
    // we need 10 bits of phase (2 for quadrant + 8 for index).
    // phase = angle * 256*4 / (2*pi) = angle * 512/pi
    //
    // Even simpler: divide the angle space into 1024 steps.
    // phase[9:0] = (angle / (2*pi)) * 1024
    //
    // For Q4.28 with range [-8,+8), 2*pi ≈ 6.283
    // We compute: phase = (angle * PHASE_SCALE) >> 28
    // where PHASE_SCALE = 2^28 * 1024 / (2*pi) = 1024 / (2*pi) * 2^28
    //                   = 162.97... * 2^28 ≈ 43,741,844,462
    // That overflows 32 bits, so we use a different approach.
    //
    // Practical approach: extract phase from angle directly.
    // 2*pi in Q4.28 = 0x6487_ED51. We need (angle mod 2*pi) / (2*pi) * 1024.
    // Since we want to avoid division, we use bit manipulation:
    //
    // angle_pos = angle mod 2*pi (reduced to [0, 2*pi))
    // We know 2*pi ≈ 6.283, which fits in 3 integer bits of Q4.28.
    // A 10-bit phase index covering [0, 2*pi) means each step = 2*pi/1024.
    // 2*pi/1024 in Q4.28 = 0x6487_ED51 >> 10 = 0x19220 (approx)
    //
    // Alternative: multiply angle by reciprocal of 2*pi to get [0,1) fraction,
    // then take upper 10 bits as phase index.
    // 1/(2*pi) in Q4.28 = 0.15915... * 2^28 = 42,722,829 = 0x028B_E60D

    localparam signed [WIDTH-1:0] RECIP_TWO_PI = 32'sh028B_E60D;  // 1/(2*pi) in Q4.28

    reg [1:0]  quadrant_r;
    reg [7:0]  table_idx_r;
    reg        negate_r;
    reg        mirror_r;

    // Intermediate: multiply angle by 1/(2*pi) to get fractional turns
    // Result is Q4.28 representing fraction of full circle
    // We only need the fractional part (lower 28 bits) → 10 upper frac bits = phase
    wire signed [63:0] phase_product = angle * RECIP_TWO_PI;
    // phase_product is Q8.56. The fractional turn is in bits [55:0].
    // We want 10 bits of phase from the fractional part.
    // Bits [55:46] of product = upper 10 bits of fractional turn
    wire [9:0] phase_raw = phase_product[55:46];

    always @(posedge clk) begin
        quadrant_r <= phase_raw[9:8];
        // Mirror index in quadrants 1 and 3
        mirror_r   <= phase_raw[8];
        if (phase_raw[8])
            table_idx_r <= ~phase_raw[7:0];  // 255 - idx
        else
            table_idx_r <= phase_raw[7:0];
        // Negate in quadrants 2 and 3
        negate_r <= phase_raw[9];
    end

    // =========================================================
    // Stage 2: Table lookup and sign application
    // =========================================================
    wire signed [WIDTH-1:0] table_val = sine_table[table_idx_r];

    always @(posedge clk) begin
        if (negate_r)
            result <= -table_val;
        else
            result <= table_val;
    end

endmodule
